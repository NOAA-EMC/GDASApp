netcdf rads_adt_j2_2018105.tmp {
dimensions:
	time = UNLIMITED ; // (11 currently)
variables:
	int adt_egm2008(time) ;
		adt_egm2008:_FillValue = 2147483647 ;
		adt_egm2008:long_name = "absolute dynamic topography (EGM2008)" ;
		adt_egm2008:standard_name = "absolute_dynamic_topography_egm2008" ;
		adt_egm2008:units = "m" ;
		adt_egm2008:scale_factor = 0.0001 ;
		adt_egm2008:coordinates = "lon lat" ;
	int adt_xgm2016(time) ;
		adt_xgm2016:_FillValue = 2147483647 ;
		adt_xgm2016:long_name = "absolute dynamic topography (XGM2016)" ;
		adt_xgm2016:standard_name = "absolute_dynamic_topography_xgm2016" ;
		adt_xgm2016:units = "m" ;
		adt_xgm2016:scale_factor = 0.0001 ;
		adt_xgm2016:coordinates = "lon lat" ;
	int cycle(time) ;
		cycle:_FillValue = 2147483647 ;
		cycle:long_name = "cycle number" ;
		cycle:field = 9905s ;
	int lat(time) ;
		lat:_FillValue = 2147483647 ;
		lat:long_name = "latitude" ;
		lat:standard_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:scale_factor = 1.e-06 ;
		lat:field = 201s ;
		lat:comment = "Positive latitude is North latitude, negative latitude is South latitude" ;
	int lon(time) ;
		lon:_FillValue = 2147483647 ;
		lon:long_name = "longitude" ;
		lon:standard_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:scale_factor = 1.e-06 ;
		lon:field = 301s ;
		lon:comment = "East longitude relative to Greenwich meridian" ;
	int pass(time) ;
		pass:_FillValue = 2147483647 ;
		pass:long_name = "pass number" ;
		pass:field = 9906s ;
	short sla(time) ;
		sla:_FillValue = 32767s ;
		sla:long_name = "sea level anomaly" ;
		sla:standard_name = "sea_surface_height_above_sea_level" ;
		sla:units = "m" ;
		sla:quality_flag = "swh sig0 range_rms range_numval flags swh_rms sig0_rms attitude" ;
		sla:scale_factor = 0.0001 ;
		sla:coordinates = "lon lat" ;
		sla:field = 0s ;
		sla:comment = "Sea level determined from satellite altitude - range - all altimetric corrections" ;
	double time_mjd(time) ;
		time_mjd:long_name = "Modified Julian Days" ;
		time_mjd:standard_name = "time" ;
		time_mjd:units = "days since 1858-11-17 00:00:00 UTC" ;
		time_mjd:field = 105s ;
		time_mjd:comment = "UTC time of measurement expressed in Modified Julian Days" ;

// global attributes:
		:Conventions = "CF-1.7" ;
		:title = "RADS 4 pass file" ;
		:institution = "EUMETSAT / NOAA / TU Delft" ;
		:source = "radar altimeter" ;
		:references = "RADS Data Manual, Version 4.2 or later" ;
		:featureType = "trajectory" ;
		:ellipsoid = "TOPEX" ;
		:ellipsoid_axis = 6378136.3 ;
		:ellipsoid_flattening = 0.00335281317789691 ;
		:filename = "rads_adt_j2_2018105.nc" ;
		:mission_name = "JASON-2" ;
		:mission_phase = "c" ;
		:log01 = "2019-01-11 | rads2nc --ymd=180415000000,180416000000 -C1,1000 -Sj2 -Vadt_egm2008,adt_xgm2016,sla,time_mjd,lon,lat,cycle,pass -Xxgm2016 -Xadt.xml -o/ftp/rads/adt//2018/rads_adt_j2_2018105.nc: RAW data from" ;
		:history = "Fri Jan 26 15:41:52 2024: ncks -d time,0,10 /scratch1/NCEPDEV/stmp4/Shastri.Paturi/forAndrew/gdas.20180415/00/adt/rads_adt_j2_2018105.nc rads_adt_j2_2018105.tmp.nc\n",
			"2019-01-11 12:29:39 : rads2nc --ymd=180415000000,180416000000 -C1,1000 -Sj2 -Vadt_egm2008,adt_xgm2016,sla,time_mjd,lon,lat,cycle,pass -Xxgm2016 -Xadt.xml -o/ftp/rads/adt//2018/rads_adt_j2_2018105.nc" ;
		:NCO = "netCDF Operators version 5.0.6 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco)" ;
data:

 adt_egm2008 = 4047, 3772, 3981, 4214, 3951, 4056, 3969, 3606, 3665, 1936, 
    2147 ;

 adt_xgm2016 = 2949, 2625, 2883, 3195, 3018, 3358, 3796, 4276, 4166, 2012, 
    2541 ;

 cycle = 349, 349, 349, 349, 349, 349, 349, 349, 349, 349, 349 ;

 lat = 49568520, 49526726, 49484908, 49443068, 49401205, 49359319, 49317410, 
    49275478, 49233524, 48516917, 48474568 ;

 lon = 153184533, 153231671, 153278722, 153325686, 153372563, 153419353, 
    153466058, 153512675, 153559207, 154337322, 154382346 ;

 pass = 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108 ;

 sla = 406, 322, 415, 554, 275, 428, 439, -392, -44, -679, -472 ;

 time_mjd = 58223.000006464, 58223.0000180141, 58223.000029564, 
    58223.000041114, 58223.0000526641, 58223.0000642141, 58223.0000757641, 
    58223.000087314, 58223.0000988641, 58223.000295214, 58223.000306764 ;
}
