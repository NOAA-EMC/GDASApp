netcdf adt.nc {
dimensions:
	Location = 100 ;
	nvars = 1 ;
variables:
	int Location(Location) ;
		Location:suggested_chunk_dim = 100LL ;
	float nvars(nvars) ;
		nvars:suggested_chunk_dim = 100LL ;

// global attributes:
		string :_ioda_layout = "ObsGroup" ;
		:_ioda_layout_version = 0 ;
		:nrecs = 1 ;
		:nvars = 1 ;
		:odb_version = 1LL ;
		:date_time = 2018041512 ;
		:nlocs = 100LL ;
		:nobs = 100LL ;
		:history = "Fri Apr 19 08:49:14 2019: ncks -d nlocs,1,50000,500 adt.orig.nc -O adt.nc" ;
		:NCO = "4.7.2" ;
data:

 Location = 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
    0, 0, 0, 0, 0, 0 ;

 nvars = 0 ;

group: MetaData {
  variables:
  	int64 dateTime(Location) ;
  		dateTime:_FillValue = -3732782400LL ;
  		string dateTime:units = "seconds since 2018-04-15T12:00:00Z" ;
  	string date_time(Location) ;
  		string date_time:_FillValue = "" ;
  	float latitude(Location) ;
  		latitude:_FillValue = 9.96921e+36f ;
  	float longitude(Location) ;
  		longitude:_FillValue = 9.96921e+36f ;
  	int sequenceNumber(Location) ;
  		sequenceNumber:_FillValue = -2147483647 ;
  	string variable_names(nvars) ;
  		string variable_names:_FillValue = "" ;
  data:

   dateTime = 8979, 37065, -10967, -28959, -42772, -24069, 28606, -17781,
      -32611, -31290, -13898, 8063, 17625, -23561, -39430, 22905, -18300,
      -31232, -23225, -38636, -18325, 8982, -9841, 29332, -10620, 37498,
      -1034, -23078, 14219, 14162, -21629, 36344, 23195, 31771, 10339, 17833,
      35703, -4052, -11549, 31202, 37231, 31403, 16181, 28642, 9593, -20577,
      8497, -3110, 17245, -39683, -24561, 8748, 23777, 5879, 17078, 600,
      -21240, -21317, 41680, -32855, 29360, -41747, -12723, -18522, 7056,
      -31791, -28776, -38385, -39168, -16351, 14451, 41413, 7784, -4273,
      -36889, -17518, -30412, -30331, -22444, -43044, 7602, 371, 34001,
      -10269, -36806, -43073, 8321, -11562, -11838, 42641, -30902, 16071,
      16374, -22526, -33032, -28369, -17501, -16309, 10748, 42986 ;

   latitude = -42.30449, -61.53271, -54.52587, 2.40806, -13.3181, -65.35713,
      -13.49405, -51.82866, 11.22875, -51.14191, 65.89512, 1.492048,
      -28.5202, -58.87149, 14.84761, -59.58656, -28.63931, -53.45946,
      -45.69531, -23.91795, -27.42865, -42.44091, -50.2743, -47.36231,
      -64.71016, -45.25023, 46.92305, -39.15643, 30.07972, 32.76525,
      30.69972, -57.81081, -65.82172, 3.266878, -52.58415, -18.54302,
      -30.36827, -60.3972, -28.85406, -24.43554, -56.09284, -14.73257,
      -60.25863, -15.23002, -64.27747, 66.14738, -19.70168, -50.90127,
      -45.91634, 27.03309, -50.4441, -31.67368, -54.68562, 53.79114,
      -52.86835, 36.03845, 48.28653, 44.95198, 6.986401, 23.08882, -48.57338,
      36.24638, 28.12075, -17.97434, 48.89173, -28.65383, 11.38542,
      -35.75763, 1.995264, -40.03509, 18.95174, 19.98642, 15.14227,
      -52.50491, -52.90968, -61.13697, -62.06583, -59.66623, -8.916806,
      -26.4584, 23.91177, 46.33038, 50.50362, -64.24638, -49.51569, -27.8661,
      -11.13248, -28.27375, -14.97766, -39.31322, -63.87175, -56.55973,
      -64.89208, -12.89731, 31.52845, 30.96179, -61.62994, -38.08575,
      -34.69767, -53.99775 ;

   longitude = -3.373801, -19.74908, 95.06168, -46.61552, 4.35299, -173.69,
      -103.4871, 119.5747, 142.6289, 175.3936, -29.76636, -23.91055,
      102.6672, -117.4293, 169.591, -36.75309, 101.5004, 178.4957, -98.71407,
      -175.7098, 100.9004, -3.265874, -160.1637, -83.9273, 124.6124,
      6.571999, -136.8072, -93.49664, -63.95547, -65.41, -63.2631, -97.47237,
      -6.842985, 58.5721, 111.8786, 107.1669, -124.3838, 78.7492, 73.26094,
      47.92515, -6.949519, 51.99478, -6.666136, -102.8136, 36.91441,
      6.947506, -15.96541, 170.7399, 91.00462, 164.346, 146.2024, -10.29815,
      52.1002, -156.9272, 83.14131, -10.65498, -50.38128, -53.59933,
      -167.6185, 137.828, -82.67605, 24.96964, 50.42411, 96.70792, -49.4618,
      158.2, -43.34373, -169.5071, 174.3347, -122.4666, -58.82631, -172.6444,
      -28.94908, 63.77332, -50.14354, 137.584, -98.06361, -90.98943,
      -79.03435, -1.207335, -32.62028, -18.51745, -164.6857, 167.3599,
      -45.90093, -1.890546, -19.34283, 72.9696, 67.16569, -147.3289,
      -155.184, -14.87442, 12.47116, -80.52476, 133.6994, -34.77795,
      139.1339, -121.1142, 127.6422, -132.5225 ;

   sequenceNumber = 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
      1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
      1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
      1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
      1, 1, 1, 1, 1, 1, 1, 1, 1 ;

   variable_names = "absolute_dynamic_topography" ;
  } // group MetaData

group: ObsError {
  variables:
  	float absoluteDynamicTopography(Location) ;
  		absoluteDynamicTopography:_FillValue = 9.96921e+36f ;
  data:

   absoluteDynamicTopography = 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1,
      0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1,
      0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1,
      0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1,
      0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1,
      0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1,
      0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1,
      0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1 ;
  } // group ObsError

group: ObsValue {
  variables:
  	float absoluteDynamicTopography(Location) ;
  		absoluteDynamicTopography:_FillValue = 9.96921e+36f ;
  data:

   absoluteDynamicTopography = 0.2886, -1.3556, -0.5692, 0.5597, 0.3317,
      -0.9281, 0.646, -0.3841, 1.1805, 0.2265, -0.3182, 0.5563, 1.1411,
      -0.4136, 1.2235, -1.1775, 0.8149, -0.0451, 0.4549, 1.1222, 0.5479,
      0.2928, 0.6877, 0.2859, -1.2493, -0.1018, 0.4664, 0.7455, 0.7465,
      0.5585, 0.6794, -0.0422, -1.4293, 0.8899, -0.9427, 1.1056, 0.9883,
      -1.0632, 1.0919, 1.3852, -0.8461, 0.9989, -1.4867, 0.7519, -1.2997,
      -0.1713, 0.5795, 0.5559, 0.3537, 1.2151, 0.2197, 0.8687, -0.7904,
      0.1346, -0.9257, 0.1562, -0.1302, -0.0695, 0.9187, 1.1942, 0.3083,
      0.2067, 0.5803, 0.8152, -0.4867, 1.291, 0.5355, 0.6636, 1.2767, 0.6614,
      0.6591, 1.3125, 0.3322, -0.6027, -0.1315, -0.9311, -0.519, -0.507,
      0.5987, 0.6005, 0.4232, 0.1729, 0.2895, -1.1387, -0.3301, 0.5248,
      0.4213, 1.0189, 0.9698, 0.6685, -1.1554, -0.942, -1.3066, 0.6466,
      1.469, 0.2632, -0.8869, 0.6544, 0.6571, -0.1728 ;
  } // group ObsValue

group: PreQc {
  variables:
  	int absoluteDynamicTopography(Location) ;
  		absoluteDynamicTopography:_FillValue = -2147483647 ;
  data:

   absoluteDynamicTopography = 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
      0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
      0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
      0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
      0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;
  } // group PreQc
}
