netcdf rads_adt_sa_2021182 {
dimensions:
	time = UNLIMITED ; // (11 currently)
variables:
	int adt_egm2008(time) ;
		adt_egm2008:_FillValue = 2147483647 ;
		adt_egm2008:long_name = "absolute dynamic topography (EGM2008)" ;
		adt_egm2008:standard_name = "absolute_dynamic_topography_egm2008" ;
		adt_egm2008:units = "m" ;
		adt_egm2008:scale_factor = 0.0001 ;
		adt_egm2008:coordinates = "lon lat" ;
	int adt_xgm2016(time) ;
		adt_xgm2016:_FillValue = 2147483647 ;
		adt_xgm2016:long_name = "absolute dynamic topography (XGM2016)" ;
		adt_xgm2016:standard_name = "absolute_dynamic_topography_xgm2016" ;
		adt_xgm2016:units = "m" ;
		adt_xgm2016:scale_factor = 0.0001 ;
		adt_xgm2016:coordinates = "lon lat" ;
	int cycle(time) ;
		cycle:_FillValue = 2147483647 ;
		cycle:long_name = "cycle number" ;
		cycle:field = 9905s ;
	int lat(time) ;
		lat:_FillValue = 2147483647 ;
		lat:long_name = "latitude" ;
		lat:standard_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:scale_factor = 1.e-06 ;
		lat:field = 201s ;
		lat:comment = "Positive latitude is North latitude, negative latitude is South latitude" ;
	int lon(time) ;
		lon:_FillValue = 2147483647 ;
		lon:long_name = "longitude" ;
		lon:standard_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:scale_factor = 1.e-06 ;
		lon:field = 301s ;
		lon:comment = "East longitude relative to Greenwich meridian" ;
	int pass(time) ;
		pass:_FillValue = 2147483647 ;
		pass:long_name = "pass number" ;
		pass:field = 9906s ;
	short sla(time) ;
		sla:_FillValue = 32767s ;
		sla:long_name = "sea level anomaly" ;
		sla:standard_name = "sea_surface_height_above_sea_level" ;
		sla:units = "m" ;
		sla:quality_flag = "swh sig0 range_rms range_numval flags peakiness" ;
		sla:scale_factor = 0.0001 ;
		sla:coordinates = "lon lat" ;
		sla:field = 0s ;
		sla:comment = "Sea level determined from satellite altitude - range - all altimetric corrections" ;
	double time_dtg(time) ;
		time_dtg:long_name = "time_dtg" ;
		time_dtg:standard_name = "time_dtg" ;
		time_dtg:units = "yyyymmddhhmmss" ;
		time_dtg:coordinates = "lon lat" ;
		time_dtg:comment = "UTC time formatted as yyyymmddhhmmss" ;
	double time_mjd(time) ;
		time_mjd:long_name = "Modified Julian Days" ;
		time_mjd:standard_name = "time" ;
		time_mjd:units = "days since 1858-11-17 00:00:00 UTC" ;
		time_mjd:field = 105s ;
		time_mjd:comment = "UTC time of measurement expressed in Modified Julian Days" ;

// global attributes:
		:Conventions = "CF-1.7" ;
		:title = "RADS 4 pass file" ;
		:institution = "EUMETSAT / NOAA / TU Delft" ;
		:source = "radar altimeter" ;
		:references = "RADS Data Manual, Version 4.2 or later" ;
		:featureType = "trajectory" ;
		:ellipsoid = "TOPEX" ;
		:ellipsoid_axis = 6378136.3 ;
		:ellipsoid_flattening = 0.00335281317789691 ;
		:filename = "rads_adt_sa_2021182.nc" ;
		:mission_name = "SARAL" ;
		:mission_phase = "b" ;
		:log01 = "2021-07-02 | /Users/rads/bin/rads2nc --ymd=20210701000000,20210702000000 -C1,1000 -Ssa -Vsla,adt_egm2008,adt_xgm2016,time_mjd,time_dtg,lon,lat,cycle,pass -X/Users/rads/cron/xgm2016 -X/Users/rads/cron/adt -X/Users/rads/cron/time_dtg -o/Users/rads/adt/2021/182/rads_adt_sa_2021182.nc: RAW data from" ;
		:history = "Mon Sep 25 17:01:33 2023: ncks -d time,0,10 rads_adt_sa_2021182.nc rads_adt_sa_2021182.ncn\n",
			"2021-07-02 21:51:14 : /Users/rads/bin/rads2nc --ymd=20210701000000,20210702000000 -C1,1000 -Ssa -Vsla,adt_egm2008,adt_xgm2016,time_mjd,time_dtg,lon,lat,cycle,pass -X/Users/rads/cron/xgm2016 -X/Users/rads/cron/adt -X/Users/rads/cron/time_dtg -o/Users/rads/adt/2021/182/rads_adt_sa_2021182.nc" ;
		:NCO = "netCDF Operators version 5.0.6 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco)" ;
data:

 adt_egm2008 = 117, 178, -117, -75, -77, -208, 157, 282, 346, 227, 424 ;

 adt_xgm2016 = -150, -98, -67, 208, 438, 374, 368, 147, 227, 206, 642 ;

 cycle = 88, 88, 88, 88, 88, 88, 88, 88, 88, 88, 88 ;

 lat = -46655742, -46594378, -46533055, -46471713, -46410368, -46349018, 
    -46287663, -46226305, -46164942, -46103576, -46042205 ;

 lon = 95661457, 95637364, 95613334, 95589341, 95565392, 95541487, 95517626, 
    95493808, 95470032, 95446300, 95422610 ;

 pass = 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63 ;

 sla = 72, 104, 84, 184, 62, -33, 108, 165, 226, 180, 238 ;

 time_dtg = 20210701000805, 20210701000806, 20210701000807, 20210701000808, 
    20210701000809, 20210701000810, 20210701000811, 20210701000812, 
    20210701000813, 20210701000814, 20210701000816 ;

 time_mjd = 59396.0056188574, 59396.0056310796, 59396.0056432929, 
    59396.005655509, 59396.0056677251, 59396.0056799412, 59396.0056921573, 
    59396.0057043734, 59396.0057165896, 59396.0057288057, 59396.0057410218 ;
}
