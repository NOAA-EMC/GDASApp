netcdf icec_mirs_snpp_2 {
dimensions:
	Scanline = 12 ;
	Field_of_view = 96 ;
	Channel = 22 ;
	Qc_dim = 4 ;
variables:
	short Atm_type(Scanline, Field_of_view) ;
		Atm_type:description = "type of atmosphere:currently missing" ;
		Atm_type:coordinates = "Longitude Latitude" ;
	short BT(Scanline, Field_of_view, Channel) ;
		BT:long_name = "Channel Temperature (K)" ;
		BT:units = "Kelvin" ;
		BT:coordinates = "Longitude Latitude Freq" ;
		BT:scale_factor = 0.01 ;
		BT:_FillValue = -999s ;
		BT:valid_range = 0, 50000 ;
	short CLW(Scanline, Field_of_view) ;
		CLW:long_name = "Cloud liquid Water (mm)" ;
		CLW:units = "mm" ;
		CLW:coordinates = "Longitude Latitude" ;
		CLW:scale_factor = 0.01 ;
		CLW:_FillValue = -999s ;
		CLW:valid_range = 0, 10000 ;
	short ChanSel(Scanline, Field_of_view, Channel) ;
		ChanSel:long_name = "Channels Selection Used in Retrieval" ;
		ChanSel:units = "1" ;
		ChanSel:coordinates = "Longitude Latitude Freq" ;
		ChanSel:_FillValue = -999s ;
		ChanSel:valid_range = 0, 1 ;
	float ChiSqr(Scanline, Field_of_view) ;
		ChiSqr:description = "Convergence rate: <3-good,>10-bad" ;
		ChiSqr:units = "1" ;
		ChiSqr:coordinates = "Longitude Latitude" ;
		ChiSqr:_FillValue = -999.f ;
		ChiSqr:valid_range = 0.f, 1000.f ;
	short CldBase(Scanline, Field_of_view) ;
		CldBase:long_name = "Cloud Base Pressure" ;
		CldBase:scale_factor = 0.1 ;
		CldBase:coordinates = "Longitude Latitude" ;
	short CldThick(Scanline, Field_of_view) ;
		CldThick:long_name = "Cloud Thickness" ;
		CldThick:scale_factor = 0.1 ;
		CldThick:coordinates = "Longitude Latitude" ;
	short CldTop(Scanline, Field_of_view) ;
		CldTop:long_name = "Cloud Top Pressure" ;
		CldTop:scale_factor = 0.1 ;
		CldTop:coordinates = "Longitude Latitude" ;
	short Emis(Scanline, Field_of_view, Channel) ;
		Emis:long_name = "Channel Emissivity" ;
		Emis:units = "1" ;
		Emis:coordinates = "Longitude Latitude Freq" ;
		Emis:scale_factor = 0.0001 ;
		Emis:_FillValue = -999s ;
		Emis:valid_range = 0, 10000 ;
	float Freq(Channel) ;
		Freq:description = "Central Frequencies (GHz)" ;
	short GWP(Scanline, Field_of_view) ;
		GWP:long_name = "Graupel Water Path (mm)" ;
		GWP:units = "mm" ;
		GWP:coordinates = "Longitude Latitude" ;
		GWP:scale_factor = 0.01 ;
		GWP:_FillValue = -999s ;
		GWP:valid_range = 0, 10000 ;
	short IWP(Scanline, Field_of_view) ;
		IWP:long_name = "Ice Water Path (mm)" ;
		IWP:units = "mm" ;
		IWP:coordinates = "Longitude Latitude" ;
		IWP:scale_factor = 0.01 ;
		IWP:_FillValue = -999s ;
		IWP:valid_range = 0, 10000 ;
	short LWP(Scanline, Field_of_view) ;
		LWP:long_name = "Liquid Water Path (mm)" ;
		LWP:units = "mm" ;
		LWP:coordinates = "Longitude Latitude" ;
		LWP:scale_factor = 0.01 ;
		LWP:_FillValue = -999s ;
		LWP:valid_range = 0, 10000 ;
	float LZ_angle(Scanline, Field_of_view) ;
		LZ_angle:long_name = "Local Zenith Angle degree" ;
		LZ_angle:units = "degrees" ;
		LZ_angle:coordinates = "Longitude Latitude" ;
		LZ_angle:_FillValue = -999.f ;
		LZ_angle:valid_range = -70.f, 70.f ;
	float Latitude(Scanline, Field_of_view) ;
		Latitude:long_name = "Latitude of the view (-90,90)" ;
		Latitude:units = "degrees" ;
		Latitude:_FillValue = -999.f ;
		Latitude:valid_range = -90.f, 90.f ;
	float Longitude(Scanline, Field_of_view) ;
		Longitude:long_name = "Longitude of the view (-180,180)" ;
		Longitude:units = "degrees" ;
		Longitude:_FillValue = -999.f ;
		Longitude:valid_range = -180.f, 180.f ;
	short Orb_mode(Scanline) ;
		Orb_mode:description = "0-ascending,1-descending" ;
		Orb_mode:units = "1" ;
		Orb_mode:_FillValue = -999s ;
		Orb_mode:valid_range = 0, 1 ;
	short Polo(Channel) ;
		Polo:description = "Polarizations" ;
	short PrecipType(Scanline, Field_of_view) ;
		PrecipType:long_name = "Precipitation Type (Frozen/Liquid)" ;
		PrecipType:coordinates = "Longitude Latitude" ;
	short Prob_SF(Scanline, Field_of_view) ;
		Prob_SF:long_name = "Probability of falling snow (%)" ;
		Prob_SF:units = "percent" ;
		Prob_SF:coordinates = "Longitude Latitude" ;
		Prob_SF:_FillValue = -999s ;
		Prob_SF:valid_range = 0, 100 ;
	short Qc(Scanline, Field_of_view, Qc_dim) ;
		Qc:description = "Qc: 0-good, 1-usable with problem, 2-bad" ;
	float RAzi_angle(Scanline, Field_of_view) ;
		RAzi_angle:long_name = "Relative Azimuth Angle 0-360 degree" ;
		RAzi_angle:coordinates = "Longitude Latitude" ;
	short RFlag(Scanline, Field_of_view) ;
		RFlag:long_name = "Rain Flag" ;
		RFlag:coordinates = "Longitude Latitude" ;
	short RR(Scanline, Field_of_view) ;
		RR:long_name = "Rain Rate (mm/hr)" ;
		RR:units = "mm/hr" ;
		RR:coordinates = "Longitude Latitude" ;
		RR:scale_factor = 0.1 ;
		RR:_FillValue = -999s ;
		RR:valid_range = 0, 1000 ;
	short RWP(Scanline, Field_of_view) ;
		RWP:long_name = "Rain Water Path (mm)" ;
		RWP:units = "mm" ;
		RWP:coordinates = "Longitude Latitude" ;
		RWP:scale_factor = 0.01 ;
		RWP:_FillValue = -999s ;
		RWP:valid_range = 0, 10000 ;
	short SFR(Scanline, Field_of_view) ;
		SFR:long_name = "Snow Fall Rate in mm/hr" ;
		SFR:units = "mm/hr" ;
		SFR:coordinates = "Longitude Latitude" ;
		SFR:scale_factor = 0.01 ;
		SFR:_FillValue = -999s ;
		SFR:valid_range = 0, 10000 ;
	short SIce(Scanline, Field_of_view) ;
		SIce:long_name = "Sea Ice Concentration (%)" ;
		SIce:units = "percent" ;
		SIce:coordinates = "Longitude Latitude" ;
		SIce:_FillValue = -999s ;
		SIce:valid_range = 0, 100 ;
	short SIce_FY(Scanline, Field_of_view) ;
		SIce_FY:long_name = "First-Year Sea Ice Concentration (%)" ;
		SIce_FY:units = "percent" ;
		SIce_FY:coordinates = "Longitude Latitude" ;
		SIce_FY:_FillValue = -999s ;
		SIce_FY:valid_range = 0, 100 ;
	short SIce_MY(Scanline, Field_of_view) ;
		SIce_MY:long_name = "Multi-Year Sea Ice Concentration (%)" ;
		SIce_MY:units = "percent" ;
		SIce_MY:coordinates = "Longitude Latitude" ;
		SIce_MY:_FillValue = -999s ;
		SIce_MY:valid_range = 0, 100 ;
	short SWE(Scanline, Field_of_view) ;
		SWE:long_name = "Snow Water Equivalent (cm)" ;
		SWE:units = "cm" ;
		SWE:coordinates = "Longitude Latitude" ;
		SWE:scale_factor = 0.01 ;
		SWE:_FillValue = -999s ;
		SWE:valid_range = 0, 10000 ;
	short SWP(Scanline, Field_of_view) ;
		SWP:long_name = "Snow Water Path" ;
		SWP:units = "mm" ;
		SWP:coordinates = "Longitude Latitude" ;
		SWP:scale_factor = 0.01 ;
		SWP:_FillValue = -999s ;
		SWP:valid_range = 0, 10000 ;
	float SZ_angle(Scanline, Field_of_view) ;
		SZ_angle:long_name = "Solar Zenith Angle (-90,90) degree" ;
		SZ_angle:coordinates = "Longitude Latitude" ;
	double ScanTime_UTC(Scanline) ;
		ScanTime_UTC:long_name = "Number of seconds since 00:00:00 UTC" ;
		ScanTime_UTC:units = "seconds" ;
		ScanTime_UTC:_FillValue = -999. ;
		ScanTime_UTC:valid_range = 0., 86400. ;
	short ScanTime_dom(Scanline) ;
		ScanTime_dom:long_name = "Calendar day of the month 1-31" ;
		ScanTime_dom:units = "days" ;
		ScanTime_dom:_FillValue = -999s ;
		ScanTime_dom:valid_range = 1, 31 ;
	short ScanTime_doy(Scanline) ;
		ScanTime_doy:long_name = "julian day 1-366" ;
		ScanTime_doy:units = "days" ;
		ScanTime_doy:_FillValue = -999s ;
		ScanTime_doy:valid_range = 1, 366 ;
	short ScanTime_hour(Scanline) ;
		ScanTime_hour:long_name = "hour of the day 0-23" ;
		ScanTime_hour:units = "hours" ;
		ScanTime_hour:_FillValue = -999s ;
		ScanTime_hour:valid_range = 0, 23 ;
	short ScanTime_minute(Scanline) ;
		ScanTime_minute:long_name = "minute of the hour 0-59" ;
		ScanTime_minute:units = "minutes" ;
		ScanTime_minute:_FillValue = -999s ;
		ScanTime_minute:valid_range = 0, 59 ;
	short ScanTime_month(Scanline) ;
		ScanTime_month:long_name = "Calendar month 1-12" ;
		ScanTime_month:units = "months" ;
		ScanTime_month:_FillValue = -999s ;
		ScanTime_month:valid_range = 1, 12 ;
	short ScanTime_second(Scanline) ;
		ScanTime_second:long_name = "second of the minute 0-59" ;
		ScanTime_second:units = "seconds" ;
		ScanTime_second:_FillValue = -999s ;
		ScanTime_second:valid_range = 0, 59 ;
	short ScanTime_year(Scanline) ;
		ScanTime_year:long_name = "Calendar Year 20XX" ;
		ScanTime_year:units = "years" ;
		ScanTime_year:_FillValue = -999s ;
		ScanTime_year:valid_range = 2011, 2050 ;
	short Sfc_type(Scanline, Field_of_view) ;
		Sfc_type:description = "type of surface:0-ocean,1-sea ice,2-land,3-snow" ;
		Sfc_type:units = "1" ;
		Sfc_type:coordinates = "Longitude Latitude" ;
		Sfc_type:_FillValue = -999s ;
		Sfc_type:valid_range = 0, 3 ;
	short Snow(Scanline, Field_of_view) ;
		Snow:long_name = "Snow Cover" ;
		Snow:units = "1" ;
		Snow:coordinates = "Longitude Latitude" ;
		Snow:_FillValue = -999s ;
		Snow:valid_range = 0, 1 ;
	short SnowGS(Scanline, Field_of_view) ;
		SnowGS:long_name = "Snow Grain Size (mm)" ;
		SnowGS:units = "mm" ;
		SnowGS:coordinates = "Longitude Latitude" ;
		SnowGS:scale_factor = 0.01 ;
		SnowGS:_FillValue = -999s ;
		SnowGS:valid_range = 0, 2000 ;
	short SurfM(Scanline, Field_of_view) ;
		SurfM:long_name = "Surface Moisture" ;
		SurfM:scale_factor = 0.1 ;
		SurfM:coordinates = "Longitude Latitude" ;
	short SurfP(Scanline, Field_of_view) ;
		SurfP:long_name = "Surface Pressure (mb)" ;
		SurfP:units = "millibars" ;
		SurfP:coordinates = "Longitude Latitude" ;
		SurfP:scale_factor = 0.1 ;
		SurfP:_FillValue = -999s ;
		SurfP:valid_range = 0, 12000 ;
	short TPW(Scanline, Field_of_view) ;
		TPW:long_name = "Total Precipitable Water (mm)" ;
		TPW:units = "mm" ;
		TPW:coordinates = "Longitude Latitude" ;
		TPW:scale_factor = 0.1 ;
		TPW:_FillValue = -999s ;
		TPW:valid_range = 0, 2000 ;
	short TSkin(Scanline, Field_of_view) ;
		TSkin:long_name = "Skin Temperature (K)" ;
		TSkin:units = "Kelvin" ;
		TSkin:coordinates = "Longitude Latitude" ;
		TSkin:scale_factor = 0.01 ;
		TSkin:_FillValue = -999s ;
		TSkin:valid_range = 0, 40000 ;
	short WindDir(Scanline, Field_of_view) ;
		WindDir:long_name = "Wind Direction" ;
		WindDir:scale_factor = 0.01 ;
		WindDir:coordinates = "Longitude Latitude" ;
	short WindSp(Scanline, Field_of_view) ;
		WindSp:long_name = "Wind Speed (m/s)" ;
		WindSp:scale_factor = 0.01 ;
		WindSp:coordinates = "Longitude Latitude" ;
	short WindU(Scanline, Field_of_view) ;
		WindU:long_name = "U-direction Wind Speed (m/s)" ;
		WindU:scale_factor = 0.01 ;
		WindU:coordinates = "Longitude Latitude" ;
	short WindV(Scanline, Field_of_view) ;
		WindV:long_name = "V-direction Wind Speed (m/s)" ;
		WindV:scale_factor = 0.01 ;
		WindV:coordinates = "Longitude Latitude" ;
	short YM(Scanline, Field_of_view, Channel) ;
		YM:long_name = "Un-Corrected Channel Temperature (K)" ;
		YM:units = "Kelvin" ;
		YM:coordinates = "Longitude Latitude Freq" ;
		YM:scale_factor = 0.01 ;
		YM:_FillValue = -999s ;
		YM:valid_range = 0, 50000 ;

// global attributes:
		:missing_value = -999 ;
		:notretrievedproduct_value = -888 ;
		:noretrieval_value = -99 ;
		:cdf_version = 4. ;
		:alg_version = 4201 ;
		:dap_version = "v11r4" ;
		:Conventions = "CF-1.5" ;
		:Metadata_Conventions = "CF-1.5, Unidata Dataset Discovery v1.0" ;
		:standard_name_vocabulary = "CF Standard Name Table (version 17, 24 March 2011)" ;
		:project = "Microwave Integrated Retrieval System" ;
		:title = "MIRS IMG" ;
		:summary = "MIRS imaging products including surface emissivity, TPW, CLW, RWP, IWP, LST." ;
		:date_created = "2021-06-30T02:00:45Z" ;
		:institution = "DOC/NOAA/NESDIS/NDE > NPOESS Data Exploitation, NESDIS, NOAA, U.S. Department of Commerce" ;
		:naming_authority = "gov.noaa.nesdis.nde" ;
		:production_site = "NSOF" ;
		:production_environment = "OE" ;
		:satellite_name = "NPP" ;
		:instrument_name = "ATMS" ;
		:creator_name = "DOC/NOAA/NESDIS/STAR > MIRS TEAM, Center for Satellite Applications and Research, NESDIS, NOAA, U.S. Department of Commerce" ;
		:creator_email = "Christopher.Grassotti@noaa.gov, Quanhua.Liu@noaa.gov, Shu-yan.Liu@noaa.gov, ryan.honeyager@noaa.gov, Yong-Keun.Lee@noaa.gov " ;
		:creator_url = "http://www.star.nesdis.noaa.gov/mirs" ;
		:publisher_name = "DOC/NOAA/NESDIS/NDE > NPOESS Data Exploitation, NESDIS, NOAA, U.S. Department of Commerce" ;
		:publisher_email = "NDE_POC@noaa.gov" ;
		:publisher_url = "http://projects.osd.noaa.gov/NDE" ;
		:Metadata_Link = "NDE product-specific output file name" ;
		:references = "http://www.star.nesdis.noaa.gov/mirs/documentation.php" ;
		:history = "Mon Jul 29 20:08:00 2024: ncks NPR-MIRS-IMG_v11r4_npp_s202106300127386_e202106300128103_c202106300200370.nc icec_mirs_snpp_2.nc\nCreated by MIRS Version 11.4" ;
		:processing_level = "NOAA Level 2 data" ;
		:source = "SATMS_npp_d20210630_t0127386_e0128103_b50120_c20210630015746003377_oebc_ops.h5" ;
		:time_coverage_start = "2021-06-30T01:27:38Z" ;
		:time_coverage_end = "2021-06-30T01:28:10Z" ;
		:cdm_data_type = "Swath" ;
		:geospatial_lat_units = "degrees_north" ;
		:geospatial_lon_units = "degrees_east" ;
		:geospatial_lat_resolution = "100" ;
		:geospatial_lon_resolution = "100" ;
		:geospatial_first_scanline_first_fov_lat = 62.49f ;
		:geospatial_first_scanline_first_fov_lon = 132.83f ;
		:geospatial_first_scanline_last_fov_lat = 71.26f ;
		:geospatial_first_scanline_last_fov_lon = -170.69f ;
		:geospatial_last_scanline_first_fov_lat = 63.63f ;
		:geospatial_last_scanline_first_fov_lon = 129.95f ;
		:geospatial_last_scanline_last_fov_lat = 72.94f ;
		:geospatial_last_scanline_last_fov_lon = -170.12f ;
		:total_number_retrievals = 1152 ;
		:percentage_optimal_retrievals = 0.1458333f ;
		:percentage_suboptimal_retrievals = 0.8541667f ;
		:percentage_bad_retrievals = 0.f ;
		:start_orbit_number = 50120 ;
		:end_orbit_number = 50120 ;
		:id = "ndepgsl-op-11_2021-06-30T02:00:45Z_0000001250129361_SATMS_npp_d20210630_t0127386_e0128103_b50120_c20210630015746003377_oebc_ops.h5" ;
		:NCO = "netCDF Operators version 5.0.6 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco)" ;
data:

 Atm_type =
  -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999,
  -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999,
  -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999,
  -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999,
  -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999,
  -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999,
  -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999,
  -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999,
  -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999,
  -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999,
  -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999,
  -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999 ;

 BT =
  27991, 27959, 27957, 27279, 25886, 24165, 22766, 22291, 22179, 22549, 
    22967, 23671, 24720, 25898, 26722, 28669, 29049, 28038, 27340, 26647, 
    25603, 24428,
  28002, 27978, 27979, 27307, 26025, 24306, 22828, 22311, 22240, 22553, 
    22969, 23527, 24540, 26060, 26772, 28553, 28964, 27935, 27272, 26517, 
    25431, 24294,
  28020, 28024, 27929, 27316, 26076, 24404, 22919, 22390, 22226, 22525, 
    22983, 23440, 24652, 25844, 26732, 28490, 28769, 27757, 27107, 26325, 
    25249, 24187,
  27978, 28027, 27910, 27323, 26154, 24487, 23022, 22415, 22227, 22517, 
    22848, 23615, 24554, 25916, 26953, 28400, 28677, 27662, 26918, 26088, 
    25013, 24021,
  27933, 28017, 27863, 27401, 26274, 24576, 23062, 22457, 22244, 22531, 
    22901, 23633, 24600, 25897, 26740, 28330, 28664, 27537, 26766, 25957, 
    24893, 24000,
  27847, 27959, 27819, 27411, 26316, 24668, 23089, 22480, 22232, 22487, 
    22959, 23623, 24589, 25700, 26784, 28293, 28581, 27330, 26576, 25772, 
    24886, 23972,
  27712, 27822, 27697, 27357, 26356, 24754, 23222, 22493, 22261, 22460, 
    22898, 23482, 24583, 25753, 26699, 28115, 28240, 26979, 26278, 25505, 
    24601, 23946,
  27526, 27620, 27485, 27227, 26330, 24777, 23199, 22582, 22310, 22489, 
    22901, 23495, 24448, 25908, 26401, 27896, 27921, 26501, 25910, 25312, 
    24562, 23831,
  27301, 27378, 27313, 27065, 26264, 24801, 23330, 22595, 22282, 22523, 
    22951, 23465, 24503, 25597, 26574, 27608, 27535, 26325, 25797, 25218, 
    24658, 23993,
  27074, 27139, 26926, 26827, 26156, 24800, 23325, 22645, 22335, 22523, 
    22889, 23568, 24358, 25721, 26538, 26963, 26821, 26019, 25567, 25076, 
    24512, 23886,
  27305, 27251, 26782, 26531, 25951, 24727, 23313, 22600, 22297, 22444, 
    22837, 23455, 24387, 25606, 26806, 26413, 25490, 25308, 25139, 24772, 
    24240, 23871,
  27246, 27177, 26617, 26410, 25910, 24786, 23417, 22617, 22247, 22544, 
    22820, 23571, 24344, 25771, 26765, 25984, 24321, 24818, 24953, 24728, 
    24221, 23724,
  27294, 27221, 26676, 26512, 25967, 24830, 23437, 22587, 22316, 22421, 
    22734, 23370, 24310, 25404, 26503, 26121, 24408, 24897, 25001, 24821, 
    24347, 23737,
  27401, 27330, 26969, 26707, 26035, 24926, 23458, 22699, 22293, 22512, 
    22859, 23383, 24206, 25629, 26513, 26540, 24868, 24976, 25042, 24727, 
    24290, 23863,
  27117, 27174, 26975, 26820, 26281, 25032, 23554, 22823, 22437, 22509, 
    22860, 23451, 24231, 25638, 26472, 26804, 26219, 25672, 25346, 25008, 
    24514, 23909,
  27139, 27196, 26935, 26843, 26312, 25034, 23601, 22828, 22390, 22485, 
    22848, 23440, 24331, 25647, 26586, 26973, 26648, 25979, 25593, 25142, 
    24519, 23993,
  27069, 27125, 26885, 26799, 26326, 25110, 23636, 22874, 22437, 22476, 
    22944, 23381, 24415, 25636, 26570, 27037, 26722, 26001, 25592, 25147, 
    24478, 23851,
  26960, 27002, 26857, 26763, 26312, 25175, 23681, 22876, 22537, 22500, 
    22878, 23300, 24237, 25309, 26522, 27081, 27083, 26195, 25744, 25196, 
    24509, 23803,
  26865, 26893, 26694, 26666, 26284, 25110, 23708, 22903, 22464, 22560, 
    22849, 23434, 24256, 25432, 26336, 26973, 27278, 26432, 25847, 25212, 
    24539, 23935,
  26818, 26835, 26671, 26650, 26243, 25173, 23722, 22929, 22448, 22522, 
    22866, 23467, 24440, 25439, 26590, 26987, 27301, 26499, 25943, 25330, 
    24679, 23895,
  26791, 26831, 26754, 26732, 26289, 25160, 23730, 22924, 22536, 22520, 
    22913, 23374, 24398, 25478, 26560, 27104, 27123, 26419, 25937, 25301, 
    24648, 23982,
  26755, 26849, 26828, 26762, 26301, 25237, 23801, 23000, 22540, 22508, 
    22887, 23311, 24360, 25574, 26797, 27187, 27075, 26375, 25882, 25289, 
    24532, 23928,
  26717, 26864, 26767, 26740, 26339, 25229, 23829, 22999, 22562, 22570, 
    22914, 23425, 24374, 25614, 26599, 27227, 27109, 26426, 25878, 25313, 
    24596, 23887,
  26720, 26877, 26746, 26756, 26321, 25245, 23836, 23015, 22593, 22520, 
    22817, 23334, 24237, 25625, 26716, 27223, 27104, 26364, 25900, 25254, 
    24589, 23892,
  26801, 26907, 26824, 26754, 26329, 25266, 23860, 23064, 22574, 22554, 
    22882, 23427, 24259, 25411, 26780, 27255, 26979, 26375, 25822, 25293, 
    24618, 24051,
  26926, 26981, 26897, 26825, 26411, 25306, 23876, 23071, 22579, 22585, 
    22942, 23342, 24251, 25250, 26634, 27299, 27020, 26365, 25947, 25284, 
    24705, 23954,
  27030, 27079, 26940, 26773, 26391, 25348, 23932, 23126, 22603, 22605, 
    22856, 23447, 24245, 25511, 26669, 27279, 27078, 26387, 25868, 25319, 
    24609, 23933,
  27064, 27150, 26863, 26782, 26373, 25284, 23886, 23119, 22604, 22630, 
    22859, 23317, 24115, 25381, 26572, 27199, 27053, 26372, 25884, 25348, 
    24620, 24093,
  27012, 27130, 26807, 26725, 26335, 25287, 23946, 23106, 22646, 22538, 
    22869, 23371, 24259, 25258, 26273, 27125, 26929, 26288, 25826, 25260, 
    24676, 24026,
  26866, 26999, 26799, 26704, 26287, 25316, 23907, 23180, 22657, 22644, 
    22829, 23378, 24189, 25490, 26500, 27066, 26840, 26247, 25747, 25259, 
    24587, 24026,
  26615, 26761, 26678, 26658, 26283, 25255, 23953, 23161, 22607, 22647, 
    22881, 23311, 24242, 25252, 26512, 27062, 26832, 26279, 25800, 25331, 
    24637, 24001,
  26271, 26438, 26534, 26520, 26252, 25340, 24010, 23151, 22650, 22532, 
    22845, 23360, 24270, 25430, 26677, 27000, 26894, 26363, 25909, 25444, 
    24715, 24094,
  25864, 26038, 26320, 26422, 26170, 25251, 23970, 23206, 22652, 22615, 
    22867, 23348, 24191, 25621, 27124, 26885, 26727, 26272, 25908, 25480, 
    24791, 24074,
  25443, 25594, 26232, 26343, 26095, 25357, 24000, 23183, 22712, 22562, 
    22799, 23287, 24329, 25271, 26463, 26735, 26572, 26186, 25804, 25338, 
    24785, 24174,
  25048, 25190, 26137, 26287, 26097, 25252, 24003, 23215, 22722, 22626, 
    22938, 23278, 24163, 25403, 26616, 26641, 26480, 26138, 25762, 25426, 
    24821, 24135,
  24718, 24900, 25948, 26182, 26029, 25268, 24035, 23215, 22709, 22593, 
    22808, 23350, 24250, 25367, 26585, 26556, 26575, 26261, 25928, 25514, 
    24872, 24321,
  24508, 24756, 25857, 26096, 26025, 25264, 24013, 23199, 22746, 22651, 
    22832, 23409, 24341, 25234, 26346, 26471, 26710, 26354, 26072, 25625, 
    25076, 24277,
  24464, 24716, 25784, 26037, 25929, 25208, 24048, 23226, 22787, 22645, 
    22862, 23414, 24236, 25237, 26223, 26332, 26759, 26432, 26085, 25674, 
    25044, 24377,
  24548, 24735, 25816, 26069, 25984, 25263, 24014, 23245, 22746, 22626, 
    22884, 23336, 24178, 25268, 26382, 26213, 26666, 26376, 26113, 25623, 
    25044, 24526,
  24653, 24752, 25951, 26112, 26004, 25244, 24016, 23275, 22734, 22646, 
    22917, 23425, 24222, 25350, 26637, 26215, 26628, 26466, 26106, 25716, 
    25134, 24480,
  24662, 24704, 25955, 26179, 26045, 25276, 24054, 23256, 22799, 22608, 
    22829, 23406, 24232, 25267, 26707, 26236, 26709, 26393, 26071, 25660, 
    25078, 24455,
  24546, 24564, 25712, 26008, 26057, 25310, 24032, 23295, 22803, 22634, 
    22890, 23312, 24054, 25238, 26424, 25952, 26879, 26443, 26070, 25530, 
    25053, 24390,
  24368, 24386, 25368, 25848, 25985, 25339, 24054, 23272, 22790, 22631, 
    22890, 23440, 24283, 25296, 26385, 25582, 26832, 26374, 25883, 25495, 
    24836, 24337,
  24235, 24255, 25312, 25812, 25925, 25295, 24057, 23259, 22814, 22645, 
    22924, 23429, 24005, 25471, 26547, 25524, 26603, 26284, 25831, 25414, 
    24729, 24143,
  24204, 24223, 25390, 25873, 25986, 25268, 24043, 23293, 22817, 22675, 
    22904, 23340, 24088, 25499, 26343, 25579, 26587, 26175, 25733, 25264, 
    24696, 24189,
  24269, 24277, 25435, 25915, 26007, 25266, 24029, 23301, 22747, 22675, 
    22880, 23303, 24145, 25367, 26524, 25463, 26593, 26203, 25757, 25272, 
    24690, 24110,
  24350, 24355, 25470, 25878, 25985, 25274, 24055, 23261, 22765, 22668, 
    22931, 23344, 24192, 25569, 26397, 25448, 26587, 26215, 25721, 25137, 
    24645, 24153,
  24398, 24415, 25455, 25929, 25994, 25299, 24053, 23266, 22813, 22697, 
    22894, 23471, 24246, 25467, 26679, 25449, 26545, 26145, 25729, 25256, 
    24535, 23965,
  24406, 24456, 25418, 25874, 25948, 25259, 24018, 23283, 22836, 22689, 
    23001, 23367, 24230, 25370, 26968, 25399, 26356, 26042, 25671, 25228, 
    24675, 24030,
  24702, 24645, 25757, 26012, 26001, 25214, 23999, 23192, 22735, 22690, 
    22851, 23377, 24137, 25338, 26615, 25585, 26339, 25837, 25450, 25088, 
    24487, 24030,
  24441, 24531, 25434, 25862, 25953, 25318, 24076, 23295, 22830, 22665, 
    22937, 23334, 24294, 25578, 26599, 25501, 26479, 26185, 25685, 25140, 
    24592, 24083,
  24466, 24553, 25510, 25892, 26011, 25262, 24026, 23295, 22808, 22677, 
    22970, 23326, 24178, 25477, 26253, 25542, 26678, 26376, 25732, 25255, 
    24629, 23984,
  24438, 24530, 25619, 25957, 26015, 25327, 24001, 23292, 22811, 22696, 
    22997, 23453, 24443, 25240, 26597, 25617, 26760, 26326, 25755, 25257, 
    24624, 24104,
  24300, 24412, 25662, 25973, 26013, 25264, 24020, 23323, 22827, 22689, 
    22886, 23410, 24240, 25304, 26691, 25620, 26804, 26451, 25855, 25322, 
    24656, 24205,
  24027, 24190, 25448, 25942, 25910, 25294, 24000, 23275, 22874, 22746, 
    23043, 23326, 24251, 25322, 26524, 25464, 26687, 26559, 26000, 25403, 
    24720, 24112,
  23597, 23826, 25229, 25700, 25908, 25276, 24009, 23285, 22885, 22678, 
    23010, 23432, 24221, 25405, 26596, 25223, 26756, 26731, 26141, 25527, 
    24733, 24105,
  22958, 23238, 25031, 25625, 25851, 25233, 24007, 23271, 22861, 22773, 
    22979, 23379, 24152, 25284, 26507, 25090, 26949, 26837, 26257, 25573, 
    24726, 24178,
  22026, 22324, 24917, 25484, 25841, 25191, 24025, 23268, 22868, 22699, 
    22962, 23400, 24291, 25312, 26701, 24865, 27088, 26885, 26263, 25654, 
    24879, 24126,
  20757, 21089, 24206, 25097, 25657, 25179, 23947, 23248, 22874, 22722, 
    22987, 23401, 24376, 25559, 26473, 23921, 26531, 26797, 26244, 25590, 
    24893, 24146,
  19255, 19651, 22840, 24226, 25277, 25067, 24004, 23278, 22852, 22832, 
    22976, 23393, 24267, 25397, 26678, 22312, 25480, 26722, 26312, 25674, 
    24881, 24220,
  17806, 18266, 21832, 23590, 25020, 24969, 23939, 23282, 22824, 22744, 
    23050, 23447, 24404, 25409, 26513, 21238, 25076, 26698, 26322, 25759, 
    25049, 24281,
  16728, 17224, 21610, 23458, 24937, 24987, 23963, 23270, 22893, 22763, 
    23079, 23399, 24310, 25493, 27029, 21326, 25254, 26760, 26407, 25867, 
    25057, 24356,
  16244, 16738, 21697, 23499, 24966, 24921, 23923, 23304, 22902, 22787, 
    23015, 23351, 24361, 25390, 26559, 21579, 25392, 26715, 26463, 25893, 
    25191, 24386,
  16398, 16854, 21683, 23549, 24957, 24973, 23919, 23236, 22870, 22898, 
    23004, 23397, 24404, 25634, 26641, 21502, 25137, 26713, 26443, 26005, 
    25167, 24454,
  17051, 17457, 21868, 23645, 24985, 24971, 23906, 23287, 22929, 22888, 
    23119, 23541, 24321, 25581, 26607, 21509, 24912, 26640, 26415, 25942, 
    25257, 24415,
  17970, 18318, 22376, 23964, 25086, 24917, 23906, 23254, 22889, 22887, 
    23000, 23466, 24270, 25532, 26557, 21959, 25061, 26682, 26515, 26029, 
    25225, 24523,
  18920, 19213, 22983, 24302, 25191, 24898, 23873, 23229, 22870, 22826, 
    23133, 23450, 24409, 25443, 26563, 22702, 25477, 26726, 26471, 26015, 
    25239, 24569,
  19704, 19977, 23372, 24532, 25290, 24911, 23853, 23256, 22901, 22837, 
    23145, 23487, 24314, 25601, 26609, 23209, 25558, 26721, 26478, 26024, 
    25367, 24559,
  20223, 20521, 23470, 24544, 25316, 24944, 23881, 23231, 22961, 22892, 
    23136, 23472, 24328, 25716, 26722, 23389, 25592, 26716, 26483, 25971, 
    25336, 24640,
  20473, 20817, 23487, 24599, 25284, 24882, 23806, 23235, 22960, 22878, 
    23097, 23471, 24394, 25701, 26801, 23329, 25647, 26712, 26411, 26018, 
    25254, 24534,
  20493, 20884, 23350, 24526, 25276, 24862, 23810, 23215, 22926, 22905, 
    23116, 23533, 24355, 25567, 26795, 23162, 25613, 26709, 26391, 25907, 
    25276, 24715,
  20344, 20759, 23345, 24569, 25241, 24844, 23798, 23244, 22936, 22835, 
    23117, 23519, 24499, 25485, 26584, 23078, 25505, 26635, 26372, 25868, 
    25207, 24573,
  20063, 20481, 23422, 24574, 25263, 24821, 23779, 23190, 22917, 22911, 
    23036, 23513, 24383, 25581, 26547, 23106, 25509, 26632, 26370, 25826, 
    25235, 24615,
  19674, 20075, 23256, 24521, 25233, 24743, 23734, 23188, 22927, 22893, 
    23048, 23452, 24389, 25629, 26791, 22968, 25600, 26608, 26376, 25787, 
    25204, 24569,
  19162, 19561, 23104, 24397, 25217, 24752, 23730, 23181, 22917, 22874, 
    23046, 23582, 24366, 25748, 26385, 22721, 25356, 26541, 26232, 25758, 
    25154, 24637,
  18534, 18924, 22785, 24295, 25147, 24697, 23706, 23176, 22956, 22960, 
    23113, 23573, 24351, 25640, 26793, 22435, 25405, 26554, 26232, 25796, 
    25111, 24485,
  17799, 18176, 22507, 24148, 25110, 24704, 23664, 23137, 22925, 22918, 
    23183, 23513, 24230, 25709, 26612, 22095, 25382, 26572, 26273, 25786, 
    25157, 24718,
  17047, 17383, 22098, 23942, 25017, 24617, 23679, 23173, 22946, 22894, 
    23107, 23470, 24475, 25674, 26644, 21755, 25264, 26585, 26312, 25863, 
    25291, 24693,
  16411, 16718, 21973, 23865, 25021, 24648, 23654, 23167, 22924, 22895, 
    23117, 23594, 24342, 25800, 26704, 21489, 25214, 26611, 26328, 25859, 
    25313, 24734,
  16121, 16394, 22072, 23908, 25019, 24640, 23666, 23132, 22994, 22982, 
    23138, 23451, 24500, 25668, 26794, 21515, 25429, 26613, 26315, 25873, 
    25251, 24608,
  16359, 16634, 22194, 23970, 25046, 24599, 23609, 23144, 22951, 22968, 
    23083, 23634, 24510, 25935, 26722, 21767, 25649, 26553, 26250, 25800, 
    25113, 24476,
  17239, 17499, 22587, 24158, 25047, 24527, 23594, 23189, 22986, 22937, 
    23153, 23601, 24591, 25868, 26847, 22215, 26024, 26500, 26156, 25685, 
    25018, 24464,
  18638, 18863, 23244, 24578, 25162, 24520, 23582, 23146, 22963, 23055, 
    23045, 23586, 24447, 25991, 27085, 22962, 26044, 26472, 26046, 25599, 
    25062, 24372,
  20218, 20382, 24161, 25035, 25267, 24526, 23566, 23131, 22998, 22978, 
    23204, 23591, 24384, 25728, 26857, 23876, 26191, 26420, 26026, 25610, 
    25045, 24333,
  21540, 21670, 24691, 25287, 25319, 24475, 23529, 23150, 23008, 22967, 
    23177, 23632, 24543, 25861, 26903, 24484, 26347, 26403, 26012, 25524, 
    24987, 24467,
  22361, 22479, 24834, 25360, 25326, 24477, 23499, 23157, 23010, 22994, 
    23170, 23676, 24728, 25788, 26895, 24436, 26268, 26410, 26032, 25574, 
    24956, 24402,
  22713, 22842, 24890, 25403, 25328, 24451, 23492, 23144, 22970, 23010, 
    23154, 23679, 24714, 25710, 26738, 24260, 26226, 26418, 26051, 25565, 
    25122, 24416,
  22851, 22984, 24907, 25370, 25287, 24371, 23448, 23146, 23030, 23000, 
    23211, 23592, 24644, 25915, 27131, 24137, 26204, 26353, 26029, 25509, 
    24971, 24363,
  23008, 23123, 25102, 25499, 25309, 24377, 23417, 23091, 23042, 22926, 
    23192, 23776, 24514, 25969, 26807, 24492, 26313, 26342, 25874, 25522, 
    24920, 24336,
  23222, 23326, 25499, 25684, 25303, 24311, 23378, 23134, 23044, 23023, 
    23190, 23743, 24872, 26050, 26601, 25317, 26794, 26360, 25935, 25492, 
    24928, 24290,
  23367, 23488, 25547, 25704, 25244, 24228, 23321, 23051, 22995, 23008, 
    23184, 23785, 24869, 25840, 26900, 25434, 26847, 26352, 25900, 25489, 
    24847, 24178,
  23323, 23485, 25463, 25672, 25172, 24193, 23299, 23088, 23035, 23083, 
    23262, 23761, 24821, 25974, 27287, 25036, 26438, 26347, 25937, 25493, 
    24907, 24260,
  23014, 23167, 25453, 25553, 25106, 24170, 23314, 23074, 23025, 23115, 
    23318, 23862, 24923, 26261, 27068, 24666, 26412, 26282, 25928, 25446, 
    24851, 24203,
  22474, 22500, 25233, 25510, 25031, 24037, 23269, 23096, 23025, 23039, 
    23339, 23892, 24857, 26390, 27096, 24035, 26320, 26301, 25915, 25450, 
    24848, 24307,
  21845, 21705, 25307, 25477, 24991, 24030, 23241, 23021, 23011, 23083, 
    23320, 23795, 24879, 26112, 26939, 23887, 26436, 26303, 25863, 25433, 
    24818, 24190,
  21569, 21335, 25420, 25499, 24851, 23912, 23219, 23037, 23000, 23107, 
    23224, 23986, 24922, 26304, 27019, 24062, 26420, 26099, 25698, 25186, 
    24584, 24025,
  27955, 27945, 27992, 27221, 25893, 24175, 22742, 22272, 22182, 22540, 
    23023, 23711, 24735, 25854, 26691, 28693, 28981, 27979, 27319, 26527, 
    25426, 24312,
  27965, 27962, 28004, 27272, 25997, 24325, 22835, 22327, 22229, 22499, 
    22990, 23742, 24696, 25878, 26560, 28598, 28953, 27896, 27198, 26354, 
    25224, 24279,
  27977, 28006, 27875, 27353, 26120, 24419, 22912, 22342, 22250, 22522, 
    22896, 23680, 24658, 26068, 26754, 28437, 28609, 27633, 26881, 26069, 
    25009, 24059,
  27924, 28001, 27887, 27351, 26121, 24510, 23026, 22411, 22239, 22557, 
    22943, 23715, 24737, 25816, 26784, 28341, 28498, 27414, 26672, 25881, 
    24812, 23779,
  27864, 27973, 27828, 27351, 26161, 24594, 23055, 22467, 22244, 22511, 
    22962, 23585, 24510, 25881, 27075, 28346, 28460, 27268, 26438, 25732, 
    24660, 23971,
  27767, 27885, 27735, 27375, 26250, 24653, 23131, 22505, 22279, 22568, 
    22909, 23568, 24572, 25910, 26593, 28245, 28253, 26910, 26239, 25540, 
    24692, 23984,
  27623, 27714, 27485, 27222, 26228, 24689, 23157, 22559, 22247, 22520, 
    22896, 23495, 24431, 25588, 26700, 27979, 27875, 26566, 25872, 25199, 
    24495, 23731,
  27423, 27480, 27321, 27033, 26192, 24743, 23237, 22565, 22302, 22471, 
    22936, 23538, 24513, 25663, 26571, 27628, 27301, 26154, 25650, 25112, 
    24400, 23797,
  27177, 27209, 27038, 26806, 26149, 24744, 23341, 22632, 22312, 22451, 
    22793, 23531, 24469, 25755, 26676, 27046, 26909, 26015, 25564, 25080, 
    24445, 23750,
  27329, 27250, 26829, 26544, 25882, 24732, 23307, 22543, 22257, 22419, 
    22754, 23374, 24336, 25421, 26632, 26476, 25225, 25098, 25052, 24801, 
    24205, 23683,
  27158, 27052, 26504, 26328, 25810, 24689, 23320, 22589, 22280, 22447, 
    22896, 23399, 24338, 25481, 26182, 25857, 24062, 24630, 24817, 24620, 
    24160, 23616,
  27110, 27006, 26439, 26298, 25837, 24779, 23431, 22633, 22268, 22472, 
    22898, 23462, 24372, 25541, 26654, 25701, 23603, 24528, 24782, 24645, 
    24103, 23675,
  27176, 27107, 26665, 26484, 25937, 24866, 23476, 22642, 22265, 22426, 
    22887, 23391, 24355, 25654, 26576, 26171, 24603, 24953, 25003, 24812, 
    24255, 23755,
  27304, 27271, 27017, 26737, 26065, 24933, 23472, 22665, 22329, 22423, 
    22815, 23408, 24310, 25494, 26712, 26760, 25728, 25472, 25236, 24818, 
    24273, 23748,
  27046, 27149, 26931, 26798, 26265, 25023, 23599, 22807, 22423, 22520, 
    22899, 23454, 24448, 25625, 26619, 26957, 26365, 25763, 25341, 24969, 
    24433, 23867,
  27096, 27188, 26970, 26874, 26344, 25085, 23615, 22823, 22460, 22531, 
    22906, 23433, 24420, 25674, 26795, 27076, 26389, 25769, 25421, 24960, 
    24458, 23858,
  27052, 27135, 26913, 26868, 26317, 25153, 23681, 22851, 22468, 22514, 
    22868, 23505, 24268, 25607, 26617, 27140, 26624, 25841, 25449, 25033, 
    24354, 23923,
  26961, 27029, 26785, 26809, 26313, 25140, 23668, 22895, 22486, 22540, 
    22870, 23513, 24227, 25451, 26597, 27148, 26904, 26049, 25580, 25063, 
    24556, 23868,
  26874, 26923, 26760, 26709, 26303, 25168, 23733, 22928, 22509, 22531, 
    22936, 23430, 24346, 25558, 26623, 27045, 26962, 26251, 25724, 25156, 
    24548, 23907,
  26822, 26843, 26726, 26713, 26256, 25161, 23733, 22960, 22563, 22576, 
    22858, 23424, 24369, 25484, 26628, 27099, 27004, 26396, 25807, 25235, 
    24568, 23974,
  26774, 26802, 26870, 26701, 26296, 25168, 23765, 22987, 22548, 22512, 
    22780, 23355, 24381, 25429, 26687, 27160, 27037, 26417, 25850, 25231, 
    24529, 23940,
  26702, 26779, 26847, 26750, 26337, 25216, 23803, 23028, 22562, 22522, 
    22801, 23412, 24304, 25710, 27009, 27265, 27157, 26532, 25946, 25318, 
    24535, 23866,
  26626, 26760, 26812, 26707, 26343, 25240, 23823, 23039, 22601, 22588, 
    22862, 23390, 24367, 25423, 26736, 27277, 27148, 26518, 25955, 25286, 
    24542, 23865,
  26597, 26760, 26748, 26688, 26308, 25306, 23877, 23026, 22562, 22497, 
    22849, 23368, 24286, 25567, 26669, 27209, 27081, 26442, 25907, 25272, 
    24540, 23890,
  26661, 26798, 26725, 26775, 26379, 25329, 23895, 23109, 22574, 22554, 
    22812, 23374, 24334, 25476, 26632, 27263, 26919, 26303, 25824, 25222, 
    24537, 23908,
  26794, 26893, 26851, 26784, 26379, 25307, 23904, 23117, 22626, 22525, 
    22765, 23347, 24139, 25606, 26588, 27301, 26947, 26321, 25837, 25282, 
    24574, 23900,
  26928, 27009, 26859, 26754, 26368, 25286, 23883, 23077, 22593, 22558, 
    22868, 23410, 24254, 25418, 26633, 27244, 26979, 26299, 25841, 25230, 
    24617, 23878,
  26995, 27083, 26854, 26689, 26323, 25298, 23924, 23115, 22609, 22530, 
    22889, 23345, 24215, 25402, 26549, 27232, 26974, 26378, 25853, 25334, 
    24654, 23905,
  26956, 27050, 26793, 26703, 26310, 25295, 23943, 23128, 22640, 22596, 
    22808, 23356, 24265, 25498, 26683, 27200, 27100, 26379, 25903, 25339, 
    24647, 23918,
  26790, 26895, 26776, 26684, 26372, 25301, 23924, 23143, 22604, 22587, 
    22816, 23326, 24158, 25622, 26452, 27184, 27122, 26449, 25963, 25425, 
    24666, 24031,
  26504, 26639, 26644, 26605, 26302, 25313, 23943, 23140, 22654, 22607, 
    22890, 23312, 24196, 25409, 26678, 27134, 27026, 26487, 26050, 25528, 
    24812, 24079,
  26146, 26319, 26422, 26503, 26218, 25324, 23961, 23180, 22689, 22609, 
    22887, 23342, 24300, 25302, 26544, 27005, 26965, 26513, 26082, 25541, 
    24882, 24099,
  25769, 25951, 26292, 26328, 26174, 25261, 23990, 23196, 22673, 22686, 
    22905, 23485, 24290, 25311, 26488, 26879, 26903, 26474, 26117, 25572, 
    24933, 24152,
  25409, 25560, 26207, 26331, 26132, 25266, 23970, 23187, 22712, 22614, 
    22831, 23437, 24243, 25544, 26344, 26818, 26904, 26560, 26135, 25666, 
    25060, 24426,
  25076, 25211, 26124, 26232, 26087, 25260, 23996, 23199, 22702, 22604, 
    22948, 23400, 24282, 25372, 26670, 26762, 26924, 26563, 26135, 25654, 
    25027, 24373,
  24788, 24961, 26085, 26184, 26079, 25267, 24039, 23249, 22751, 22711, 
    22878, 23407, 24357, 25504, 26381, 26603, 26813, 26498, 26157, 25649, 
    25218, 24473,
  24597, 24833, 25992, 26098, 26025, 25274, 23979, 23245, 22750, 22671, 
    22901, 23335, 24314, 25304, 26500, 26457, 26656, 26344, 26032, 25604, 
    25122, 24408,
  24547, 24789, 25931, 26055, 25988, 25190, 24010, 23249, 22762, 22693, 
    22837, 23315, 24288, 25198, 26688, 26404, 26599, 26300, 26025, 25697, 
    25161, 24435,
  24604, 24792, 25904, 26078, 25976, 25223, 24014, 23235, 22761, 22675, 
    22948, 23321, 24230, 25403, 26612, 26324, 26685, 26410, 26046, 25653, 
    25090, 24477,
  24671, 24787, 25950, 26125, 26054, 25276, 24048, 23251, 22832, 22643, 
    22935, 23430, 24317, 25378, 26679, 26218, 26712, 26363, 26074, 25738, 
    25072, 24478,
  24652, 24723, 25907, 26097, 26060, 25287, 24043, 23298, 22814, 22697, 
    22956, 23356, 24373, 25379, 26516, 26164, 26716, 26332, 26010, 25646, 
    25067, 24539,
  24535, 24591, 25553, 25961, 25978, 25275, 24039, 23305, 22781, 22677, 
    22848, 23381, 24244, 25567, 26791, 25852, 26713, 26384, 25961, 25578, 
    25048, 24387,
  24399, 24463, 25329, 25821, 25946, 25308, 24072, 23300, 22811, 22628, 
    22915, 23313, 24219, 25502, 26641, 25487, 26672, 26343, 25954, 25542, 
    24985, 24415,
  24350, 24414, 25305, 25807, 25938, 25294, 24026, 23289, 22840, 22757, 
    22925, 23292, 24284, 25315, 26606, 25401, 26660, 26369, 25943, 25561, 
    25030, 24482,
  24418, 24469, 25398, 25890, 25987, 25293, 24057, 23300, 22800, 22700, 
    22951, 23442, 24209, 25345, 26288, 25461, 26650, 26311, 25893, 25499, 
    24908, 24381,
  24559, 24585, 25588, 25950, 26041, 25316, 24033, 23320, 22819, 22657, 
    22847, 23342, 24316, 25253, 26197, 25613, 26700, 26317, 25882, 25406, 
    24915, 24275,
  24662, 24685, 25832, 26056, 26070, 25304, 24062, 23281, 22868, 22659, 
    22972, 23347, 24269, 25212, 26109, 25710, 26737, 26286, 25819, 25383, 
    24730, 24238,
  24673, 24725, 25762, 26037, 26068, 25264, 24070, 23288, 22863, 22766, 
    22903, 23405, 24157, 25437, 26663, 25719, 26840, 26310, 25828, 25297, 
    24792, 24124,
  24610, 24713, 25476, 25862, 26015, 25315, 24062, 23284, 22819, 22694, 
    22965, 23372, 24248, 25289, 26600, 25501, 26681, 26294, 25797, 25343, 
    24735, 24142,
  24552, 24680, 25402, 25865, 25961, 25271, 24053, 23321, 22815, 22737, 
    22869, 23382, 24106, 25377, 26335, 25351, 26629, 26393, 25795, 25230, 
    24690, 24088,
  24541, 24652, 25407, 25912, 25998, 25303, 24073, 23308, 22845, 22774, 
    22924, 23405, 24205, 25333, 26570, 25392, 26754, 26422, 25812, 25226, 
    24613, 24135,
  24568, 24635, 25485, 25904, 26032, 25312, 24071, 23317, 22914, 22742, 
    23014, 23506, 24243, 25410, 26559, 25418, 26753, 26476, 25851, 25359, 
    24651, 24101,
  24550, 24600, 25529, 25944, 26013, 25286, 24091, 23326, 22887, 22707, 
    22995, 23365, 24231, 25435, 26688, 25474, 26779, 26491, 25943, 25442, 
    24690, 24101,
  24407, 24489, 25538, 25966, 25991, 25317, 24031, 23286, 22871, 22689, 
    22885, 23446, 24282, 25393, 26301, 25564, 26738, 26450, 25953, 25419, 
    24766, 24323,
  24121, 24280, 25468, 25895, 25986, 25261, 24021, 23312, 22883, 22717, 
    23036, 23433, 24384, 25285, 26834, 25442, 26613, 26443, 25905, 25407, 
    24728, 24130,
  23708, 23949, 25065, 25626, 25869, 25230, 24048, 23331, 22845, 22775, 
    22963, 23418, 24298, 25442, 26810, 25072, 26569, 26469, 25963, 25413, 
    24716, 24176,
  23146, 23437, 24604, 25317, 25691, 25249, 24004, 23284, 22856, 22756, 
    22977, 23474, 24254, 25356, 26440, 24597, 26259, 26569, 26073, 25484, 
    24792, 24190,
  22350, 22649, 24608, 25330, 25765, 25168, 24025, 23278, 22933, 22814, 
    23018, 23344, 24298, 25224, 26717, 24567, 26423, 26725, 26176, 25590, 
    24849, 24204,
  21229, 21563, 24695, 25384, 25742, 25156, 23989, 23288, 22919, 22702, 
    23010, 23485, 24310, 25391, 26449, 24634, 26881, 26795, 26210, 25601, 
    24920, 24365,
  19833, 20248, 23875, 24917, 25531, 25144, 23976, 23324, 22911, 22784, 
    23037, 23393, 24351, 25418, 26285, 23540, 26290, 26785, 26313, 25801, 
    24922, 24265,
  18420, 18926, 22606, 24068, 25219, 25041, 23942, 23263, 22886, 22801, 
    23063, 23445, 24296, 25414, 26525, 22045, 25278, 26682, 26434, 25881, 
    25064, 24400,
  17327, 17895, 21768, 23573, 24974, 24953, 23936, 23286, 22858, 22886, 
    23007, 23389, 24259, 25470, 26532, 21343, 25101, 26657, 26415, 25926, 
    25116, 24481,
  16825, 17410, 21737, 23555, 24936, 24903, 23912, 23301, 22920, 22844, 
    23079, 23534, 24194, 25619, 26424, 21570, 25264, 26691, 26410, 25909, 
    25168, 24431,
  16994, 17544, 22101, 23739, 24984, 24953, 23881, 23270, 22915, 22843, 
    23022, 23443, 24372, 25694, 26535, 21747, 25287, 26682, 26451, 25972, 
    25257, 24526,
  17685, 18168, 22317, 23897, 25029, 24947, 23885, 23265, 22888, 22818, 
    23052, 23445, 24315, 25551, 26690, 21958, 25151, 26638, 26396, 25951, 
    25207, 24520,
  18624, 19016, 22794, 24232, 25173, 24958, 23907, 23243, 22921, 22872, 
    23132, 23553, 24257, 25528, 26816, 22504, 25380, 26659, 26447, 25976, 
    25310, 24579,
  19533, 19844, 23343, 24465, 25238, 24897, 23856, 23254, 22898, 22876, 
    23060, 23460, 24293, 25613, 26685, 23151, 25591, 26752, 26465, 26000, 
    25254, 24586,
  20223, 20509, 23559, 24655, 25281, 24915, 23904, 23243, 22895, 22829, 
    23134, 23449, 24339, 25582, 27107, 23481, 25641, 26712, 26451, 26028, 
    25330, 24730,
  20648, 20958, 23630, 24621, 25334, 24927, 23818, 23253, 22947, 22926, 
    23098, 23531, 24519, 25558, 26497, 23464, 25675, 26700, 26429, 26100, 
    25370, 24704,
  20860, 21192, 23449, 24551, 25257, 24878, 23849, 23228, 22928, 22849, 
    23061, 23484, 24309, 25429, 26606, 23349, 25512, 26659, 26427, 26004, 
    25320, 24766,
  20917, 21251, 23495, 24563, 25334, 24852, 23762, 23229, 22947, 22916, 
    23126, 23537, 24275, 25450, 26635, 23293, 25465, 26585, 26359, 25907, 
    25240, 24633,
  20859, 21186, 23639, 24689, 25282, 24855, 23778, 23290, 22934, 22907, 
    23167, 23542, 24294, 25665, 26801, 23409, 25669, 26604, 26311, 25854, 
    25152, 24611,
  20687, 21026, 23721, 24702, 25336, 24778, 23783, 23203, 22947, 22905, 
    23106, 23549, 24395, 25687, 26962, 23521, 25604, 26603, 26275, 25787, 
    25198, 24486,
  20388, 20755, 23626, 24679, 25293, 24782, 23762, 23287, 22956, 22898, 
    23061, 23531, 24429, 25754, 26671, 23436, 25739, 26621, 26288, 25878, 
    25238, 24620,
  19926, 20334, 23501, 24640, 25264, 24765, 23744, 23224, 22964, 22890, 
    23201, 23503, 24581, 25747, 26753, 23273, 25576, 26510, 26219, 25850, 
    25214, 24661,
  19299, 19709, 23233, 24487, 25204, 24760, 23747, 23236, 22944, 22921, 
    23100, 23573, 24398, 25691, 26828, 23015, 25576, 26596, 26274, 25850, 
    25317, 24737,
  18509, 18896, 22844, 24303, 25157, 24759, 23729, 23138, 22972, 22926, 
    23173, 23635, 24485, 25551, 26328, 22620, 25583, 26600, 26268, 25915, 
    25273, 24649,
  17643, 17988, 22447, 24126, 25064, 24607, 23679, 23169, 22960, 22925, 
    23083, 23571, 24484, 25928, 27006, 22173, 25546, 26576, 26279, 25941, 
    25383, 24777,
  16856, 17189, 22168, 23945, 25074, 24633, 23629, 23171, 22998, 22955, 
    23124, 23621, 24463, 25750, 26828, 21849, 25509, 26587, 26274, 25918, 
    25366, 24758,
  16421, 16736, 22110, 23940, 25032, 24628, 23642, 23167, 22947, 22971, 
    23171, 23573, 24576, 25892, 27078, 21794, 25785, 26588, 26255, 25826, 
    25278, 24706,
  16566, 16874, 22249, 24058, 25050, 24568, 23585, 23140, 22917, 22968, 
    23175, 23713, 24525, 25738, 26747, 21959, 25812, 26509, 26106, 25737, 
    25077, 24533,
  17407, 17673, 22572, 24240, 25042, 24565, 23598, 23176, 22983, 22917, 
    23136, 23682, 24381, 25735, 26778, 22268, 25907, 26484, 26074, 25682, 
    25078, 24508,
  18792, 19007, 23352, 24596, 25132, 24502, 23593, 23133, 22970, 22949, 
    23208, 23559, 24566, 25782, 27224, 23020, 26001, 26406, 26061, 25578, 
    25065, 24449,
  20352, 20519, 24206, 25086, 25220, 24491, 23531, 23141, 23007, 22989, 
    23134, 23627, 24447, 25744, 26703, 23962, 26212, 26404, 25986, 25565, 
    24983, 24464,
  21648, 21801, 24769, 25326, 25307, 24457, 23498, 23146, 23000, 22969, 
    23184, 23736, 24722, 25768, 26869, 24550, 26350, 26430, 26035, 25615, 
    25035, 24599,
  22449, 22590, 24907, 25418, 25285, 24440, 23468, 23120, 23002, 22977, 
    23174, 23689, 24746, 25869, 26929, 24525, 26276, 26387, 26054, 25646, 
    25154, 24433,
  22783, 22912, 24930, 25389, 25295, 24405, 23436, 23130, 22971, 22998, 
    23178, 23801, 24680, 25968, 27054, 24428, 26216, 26467, 26087, 25650, 
    25099, 24580,
  22888, 22999, 24973, 25404, 25240, 24381, 23448, 23141, 23022, 23037, 
    23264, 23684, 24541, 25915, 27122, 24313, 26206, 26380, 25969, 25569, 
    25011, 24514,
  22992, 23085, 24983, 25439, 25236, 24334, 23387, 23066, 22996, 23026, 
    23185, 23865, 24766, 26000, 27006, 24436, 26241, 26340, 25957, 25657, 
    25037, 24441,
  23163, 23259, 25192, 25522, 25238, 24276, 23378, 23062, 22986, 23028, 
    23251, 23654, 24809, 25962, 27007, 24881, 26441, 26250, 25828, 25472, 
    24822, 24334,
  23321, 23444, 25322, 25579, 25174, 24247, 23290, 23073, 23045, 23014, 
    23191, 23712, 24764, 26090, 27147, 24914, 26432, 26228, 25901, 25462, 
    24894, 24415,
  23368, 23526, 25278, 25550, 25129, 24164, 23299, 23093, 22974, 23007, 
    23249, 23802, 24650, 25991, 27217, 24656, 26215, 26216, 25829, 25460, 
    24882, 24271,
  23199, 23336, 25346, 25579, 25090, 24108, 23318, 23088, 23025, 23041, 
    23299, 23765, 24783, 26229, 26996, 24576, 26309, 26194, 25833, 25357, 
    24878, 24287,
  22793, 22802, 25399, 25560, 24978, 24061, 23227, 23060, 23023, 23053, 
    23241, 23889, 24902, 26209, 26917, 24295, 26322, 26243, 25793, 25429, 
    24761, 24205,
  22249, 22106, 25388, 25571, 24992, 23990, 23220, 23078, 23009, 22982, 
    23324, 23975, 24971, 26157, 27281, 24225, 26407, 26237, 25857, 25437, 
    24821, 24308,
  22001, 21771, 25490, 25501, 24931, 23912, 23153, 23036, 23054, 23109, 
    23342, 23926, 24888, 26179, 27247, 24237, 26335, 26197, 25726, 25296, 
    24707, 24023,
  27898, 27874, 27938, 27280, 25917, 24180, 22764, 22262, 22240, 22528, 
    22965, 23760, 24848, 25985, 26602, 28738, 28901, 27713, 27066, 26349, 
    25228, 24119,
  27905, 27892, 27934, 27309, 25959, 24318, 22829, 22315, 22202, 22550, 
    22981, 23550, 24634, 25844, 26816, 28569, 28729, 27573, 26820, 26064, 
    24999, 23952,
  27908, 27935, 27791, 27247, 26054, 24410, 22940, 22348, 22249, 22495, 
    22966, 23666, 24714, 25715, 26629, 28434, 28416, 27279, 26484, 25747, 
    24728, 23800,
  27845, 27930, 27803, 27276, 26179, 24501, 23003, 22437, 22255, 22556, 
    22993, 23562, 24607, 25843, 26821, 28259, 28244, 27090, 26273, 25554, 
    24607, 23732,
  27779, 27888, 27679, 27265, 26165, 24560, 23049, 22434, 22255, 22538, 
    22976, 23439, 24551, 25832, 26589, 28223, 28038, 26807, 26006, 25460, 
    24568, 23898,
  27680, 27771, 27575, 27221, 26119, 24622, 23117, 22455, 22214, 22473, 
    22903, 23642, 24503, 25782, 26622, 28026, 27706, 26406, 25792, 25200, 
    24525, 23817,
  27532, 27567, 27374, 27094, 26182, 24657, 23175, 22538, 22322, 22543, 
    22873, 23503, 24487, 25847, 26904, 27726, 27396, 26207, 25626, 25082, 
    24436, 23792,
  27323, 27313, 27125, 26875, 26084, 24684, 23228, 22576, 22295, 22531, 
    22910, 23549, 24424, 25999, 26827, 27234, 26847, 26018, 25583, 25088, 
    24462, 23830,
  27468, 27361, 26842, 26535, 25850, 24667, 23262, 22501, 22268, 22573, 
    22861, 23435, 24513, 25807, 26696, 26607, 25978, 25603, 25315, 24915, 
    24293, 23757,
  27209, 27083, 26447, 26265, 25772, 24681, 23293, 22545, 22268, 22463, 
    22898, 23473, 24385, 25604, 26703, 25924, 24057, 24594, 24784, 24653, 
    24235, 23816,
  27041, 26897, 26403, 26176, 25751, 24717, 23377, 22589, 22311, 22457, 
    22890, 23496, 24485, 25495, 26774, 25659, 24287, 24896, 24963, 24696, 
    24216, 23730,
  27007, 26874, 26501, 26276, 25818, 24784, 23411, 22610, 22308, 22483, 
    22898, 23526, 24391, 25567, 26490, 25941, 24311, 24810, 24893, 24640, 
    24196, 23723,
  27086, 27008, 26657, 26540, 25978, 24876, 23445, 22680, 22302, 22477, 
    22997, 23376, 24386, 25472, 26698, 26472, 25349, 25271, 25128, 24789, 
    24285, 23922,
  26845, 26943, 26787, 26715, 26138, 24951, 23528, 22798, 22420, 22559, 
    22887, 23391, 24449, 25644, 26313, 26801, 26374, 25830, 25401, 24960, 
    24410, 23852,
  26980, 27101, 26854, 26751, 26187, 25000, 23537, 22839, 22434, 22539, 
    22918, 23420, 24371, 25438, 26656, 26997, 26415, 25685, 25308, 24846, 
    24349, 23881,
  27053, 27159, 26906, 26800, 26268, 25043, 23598, 22867, 22466, 22536, 
    22948, 23421, 24239, 25561, 26658, 27120, 26184, 25632, 25278, 24923, 
    24342, 23812,
  27034, 27132, 26926, 26781, 26332, 25063, 23633, 22878, 22503, 22522, 
    22915, 23451, 24423, 25704, 26591, 27156, 26550, 25828, 25430, 24984, 
    24536, 23903,
  26958, 27053, 26832, 26772, 26231, 25171, 23637, 22901, 22531, 22600, 
    22895, 23486, 24254, 25484, 26812, 27156, 26774, 26013, 25574, 25071, 
    24453, 23875,
  26867, 26953, 26739, 26712, 26284, 25148, 23689, 22972, 22517, 22562, 
    22815, 23417, 24241, 25672, 26636, 27117, 26807, 26215, 25663, 25126, 
    24534, 23947,
  26792, 26847, 26810, 26750, 26251, 25169, 23758, 22983, 22541, 22675, 
    22878, 23420, 24440, 25600, 26794, 27109, 27012, 26281, 25766, 25218, 
    24528, 23921,
  26708, 26750, 26801, 26724, 26288, 25201, 23794, 23008, 22515, 22588, 
    22948, 23418, 24393, 25620, 26755, 27179, 27100, 26476, 25954, 25313, 
    24654, 23954,
  26602, 26666, 26747, 26682, 26287, 25154, 23789, 23007, 22581, 22572, 
    22954, 23421, 24301, 25644, 26826, 27203, 27096, 26510, 25975, 25488, 
    24629, 23914,
  26495, 26601, 26675, 26679, 26298, 25181, 23817, 23003, 22621, 22615, 
    22843, 23368, 24270, 25546, 26499, 27182, 27099, 26484, 25922, 25362, 
    24590, 23979,
  26442, 26584, 26628, 26684, 26303, 25261, 23836, 23046, 22590, 22662, 
    22929, 23404, 24171, 25739, 26490, 27206, 27144, 26508, 25957, 25354, 
    24615, 23904,
  26492, 26633, 26739, 26709, 26306, 25250, 23875, 23071, 22629, 22628, 
    22987, 23413, 24442, 25484, 26633, 27240, 27212, 26540, 26066, 25373, 
    24670, 23954,
  26630, 26751, 26791, 26782, 26321, 25273, 23894, 23090, 22618, 22593, 
    22925, 23396, 24217, 25388, 26551, 27298, 27172, 26581, 26053, 25383, 
    24642, 24040,
  26790, 26886, 26833, 26685, 26340, 25255, 23932, 23109, 22635, 22635, 
    22931, 23428, 24259, 25450, 26741, 27191, 27062, 26537, 26056, 25462, 
    24754, 23972,
  26890, 26969, 26788, 26688, 26272, 25283, 23915, 23079, 22637, 22609, 
    22914, 23411, 24242, 25495, 26431, 27176, 27068, 26580, 26081, 25528, 
    24799, 24005,
  26872, 26933, 26784, 26738, 26357, 25328, 23906, 23137, 22681, 22612, 
    22921, 23349, 24283, 25508, 26373, 27219, 27244, 26610, 26111, 25577, 
    24785, 24105,
  26711, 26770, 26691, 26707, 26306, 25306, 23998, 23125, 22709, 22592, 
    22855, 23365, 24176, 25425, 26419, 27185, 27278, 26644, 26172, 25538, 
    24861, 24171,
  26427, 26510, 26629, 26612, 26283, 25293, 23979, 23181, 22700, 22594, 
    22842, 23373, 24177, 25341, 26657, 27141, 27264, 26660, 26175, 25641, 
    24975, 24321,
  26092, 26210, 26429, 26531, 26217, 25323, 24007, 23150, 22726, 22608, 
    22952, 23454, 24265, 25475, 26831, 27054, 27220, 26729, 26263, 25785, 
    25052, 24373,
  25760, 25891, 26314, 26375, 26161, 25317, 23977, 23208, 22714, 22611, 
    22879, 23336, 24353, 25223, 26501, 26906, 27097, 26625, 26249, 25765, 
    25008, 24394,
  25450, 25561, 26231, 26360, 26172, 25266, 24015, 23222, 22730, 22645, 
    22931, 23411, 24184, 25367, 26431, 26845, 26949, 26618, 26226, 25891, 
    25230, 24534,
  25152, 25257, 26146, 26326, 26117, 25248, 24007, 23212, 22748, 22617, 
    22899, 23306, 24222, 25312, 26355, 26760, 26962, 26571, 26254, 25730, 
    25217, 24554,
  24878, 25018, 26059, 26239, 26065, 25270, 24036, 23261, 22779, 22707, 
    22894, 23333, 24187, 25521, 26451, 26614, 26982, 26599, 26241, 25856, 
    25229, 24667,
  24685, 24871, 25915, 26132, 26019, 25243, 24004, 23241, 22775, 22670, 
    22918, 23366, 24262, 25337, 26518, 26432, 26744, 26417, 26165, 25761, 
    25242, 24582,
  24619, 24796, 25875, 26048, 25984, 25207, 23990, 23251, 22743, 22618, 
    22843, 23318, 24253, 25333, 26450, 26323, 26606, 26337, 25963, 25649, 
    25191, 24616,
  24649, 24772, 25810, 26013, 25957, 25226, 24036, 23270, 22769, 22631, 
    22924, 23477, 24101, 25142, 26198, 26196, 26550, 26216, 25909, 25573, 
    25101, 24544,
  24688, 24756, 25858, 26057, 25973, 25245, 23948, 23203, 22804, 22653, 
    22926, 23357, 24129, 25276, 26441, 26156, 26513, 26234, 25860, 25536, 
    25160, 24559,
  24654, 24705, 25716, 25959, 26008, 25251, 24026, 23257, 22787, 22627, 
    22890, 23285, 24226, 25379, 26924, 25968, 26610, 26334, 25929, 25592, 
    25154, 24647,
  24554, 24618, 25481, 25933, 25908, 25247, 24007, 23217, 22833, 22673, 
    22956, 23359, 24305, 25330, 26726, 25651, 26459, 26247, 25907, 25517, 
    25085, 24501,
  24476, 24570, 25438, 25895, 25993, 25271, 24031, 23241, 22804, 22693, 
    22897, 23334, 24228, 25425, 26104, 25540, 26511, 26243, 25907, 25525, 
    24983, 24543,
  24523, 24629, 25603, 25971, 25990, 25251, 24061, 23312, 22811, 22621, 
    22839, 23318, 24121, 25378, 26653, 25609, 26712, 26326, 25924, 25537, 
    25041, 24442,
  24697, 24792, 25615, 26035, 25994, 25309, 24023, 23268, 22787, 22682, 
    22889, 23401, 24144, 25332, 26332, 25653, 26768, 26391, 25991, 25500, 
    25047, 24542,
  24918, 24986, 25741, 26089, 26050, 25307, 24068, 23287, 22847, 22699, 
    22904, 23395, 24177, 25232, 26816, 25706, 26782, 26346, 25912, 25495, 
    24977, 24509,
  25053, 25122, 25974, 26171, 26099, 25292, 24035, 23322, 22824, 22727, 
    22971, 23350, 24264, 25407, 26447, 25964, 26831, 26359, 25868, 25447, 
    24907, 24433,
  25049, 25159, 25949, 26110, 26131, 25289, 24061, 23288, 22857, 22748, 
    22829, 23345, 24098, 25234, 26519, 25983, 26840, 26346, 25857, 25423, 
    24848, 24371,
  24945, 25116, 25840, 26074, 26056, 25282, 24050, 23317, 22841, 22711, 
    22976, 23395, 24316, 25172, 26375, 25800, 26794, 26359, 25840, 25357, 
    24822, 24236,
  24849, 25041, 25713, 26006, 26062, 25271, 24011, 23306, 22847, 22736, 
    22982, 23317, 24229, 25575, 26746, 25656, 26743, 26422, 25824, 25225, 
    24688, 24195,
  24818, 24974, 25691, 25992, 25984, 25289, 24007, 23316, 22879, 22701, 
    22960, 23406, 24239, 25317, 26811, 25676, 26787, 26407, 25793, 25326, 
    24771, 24175,
  24842, 24932, 25644, 25987, 26053, 25279, 24045, 23332, 22905, 22739, 
    22965, 23406, 24376, 25514, 26419, 25625, 26828, 26526, 25963, 25323, 
    24700, 24143,
  24821, 24891, 25745, 26056, 26046, 25328, 24050, 23320, 22911, 22738, 
    22985, 23385, 24349, 25551, 26860, 25639, 26812, 26536, 25986, 25356, 
    24765, 24276,
  24664, 24774, 25701, 26057, 26026, 25241, 24014, 23288, 22868, 22714, 
    22910, 23449, 24129, 25435, 26668, 25695, 26763, 26509, 25941, 25365, 
    24771, 24036,
  24357, 24548, 25537, 25943, 25964, 25264, 24056, 23271, 22871, 22711, 
    22958, 23397, 24243, 25295, 26316, 25524, 26496, 26321, 25789, 25303, 
    24644, 24211,
  23941, 24201, 25185, 25717, 25876, 25246, 23993, 23337, 22830, 22754, 
    22997, 23352, 24345, 25365, 26321, 25122, 26521, 26447, 25924, 25415, 
    24688, 24137,
  23418, 23706, 24749, 25456, 25769, 25150, 23963, 23269, 22864, 22727, 
    23011, 23494, 24150, 25347, 26619, 24577, 26446, 26591, 26074, 25485, 
    24752, 24163,
  22713, 22995, 24642, 25350, 25743, 25159, 23974, 23295, 22871, 22775, 
    23001, 23304, 24243, 25406, 26725, 24460, 26218, 26638, 26184, 25585, 
    24829, 24158,
  21715, 22033, 24735, 25378, 25711, 25211, 24042, 23294, 22898, 22782, 
    22937, 23422, 24192, 25442, 26772, 24715, 26632, 26810, 26309, 25676, 
    24900, 24292,
  20438, 20846, 24407, 25193, 25678, 25152, 24001, 23317, 22925, 22828, 
    23014, 23471, 24153, 25332, 26456, 24342, 26609, 26887, 26350, 25754, 
    25009, 24466,
  19112, 19622, 23307, 24471, 25346, 25099, 23978, 23277, 22906, 22823, 
    23048, 23312, 24438, 25338, 26288, 23023, 25976, 26776, 26374, 25846, 
    25093, 24379,
  18070, 18652, 22225, 23771, 25104, 24994, 23947, 23310, 22922, 22828, 
    22954, 23387, 24355, 25440, 26331, 21783, 25020, 26491, 26368, 25860, 
    25057, 24307,
  17600, 18204, 22074, 23639, 24997, 24929, 23906, 23322, 22899, 22800, 
    23070, 23418, 24306, 25400, 26600, 21766, 25128, 26562, 26391, 25905, 
    25128, 24311,
  17790, 18357, 22414, 23953, 25085, 24938, 23923, 23270, 22911, 22831, 
    22970, 23502, 24298, 25548, 26735, 22218, 25531, 26632, 26376, 25942, 
    25142, 24367,
  18480, 18968, 22729, 24125, 25156, 24887, 23882, 23262, 22905, 22772, 
    22995, 23365, 24183, 25481, 26026, 22529, 25475, 26654, 26404, 25954, 
    25174, 24460,
  19368, 19753, 23195, 24438, 25217, 24946, 23896, 23243, 22915, 22791, 
    22964, 23478, 24200, 25346, 26493, 22921, 25393, 26688, 26442, 26041, 
    25276, 24528,
  20175, 20476, 23695, 24741, 25354, 24964, 23857, 23271, 22897, 22814, 
    22986, 23392, 24332, 25227, 26751, 23552, 25747, 26674, 26459, 26040, 
    25303, 24594,
  20741, 21026, 23829, 24765, 25356, 24895, 23837, 23228, 22918, 22857, 
    22994, 23376, 24301, 25533, 26496, 23743, 25859, 26670, 26466, 25943, 
    25341, 24550,
  21066, 21380, 23750, 24752, 25307, 24910, 23847, 23271, 22963, 22831, 
    23023, 23372, 24355, 25313, 26816, 23629, 25743, 26657, 26389, 25971, 
    25298, 24692,
  21238, 21554, 23681, 24683, 25301, 24872, 23814, 23242, 22875, 22879, 
    23012, 23414, 24303, 25523, 26684, 23488, 25624, 26638, 26386, 25819, 
    25235, 24613,
  21310, 21593, 23791, 24745, 25321, 24897, 23771, 23237, 22955, 22901, 
    23065, 23435, 24360, 25462, 26869, 23587, 25696, 26600, 26304, 25809, 
    25137, 24501,
  21303, 21552, 23978, 24847, 25351, 24826, 23823, 23249, 22936, 22861, 
    23035, 23510, 24289, 25656, 26680, 23727, 25762, 26576, 26299, 25818, 
    25188, 24612,
  21196, 21461, 23938, 24820, 25374, 24789, 23790, 23187, 22928, 22830, 
    23119, 23518, 24356, 25610, 26796, 23786, 25728, 26551, 26297, 25751, 
    25095, 24620,
  20964, 21281, 23861, 24844, 25340, 24815, 23759, 23189, 22974, 22906, 
    23063, 23511, 24493, 25523, 26671, 23773, 25801, 26578, 26248, 25818, 
    25147, 24600,
  20563, 20943, 23706, 24701, 25282, 24756, 23714, 23171, 22975, 22881, 
    23090, 23544, 24425, 25532, 26803, 23660, 25993, 26582, 26193, 25795, 
    25200, 24648,
  19980, 20372, 23580, 24632, 25224, 24720, 23689, 23176, 22938, 22879, 
    23119, 23479, 24466, 25678, 27173, 23491, 25887, 26610, 26262, 25926, 
    25353, 24731,
  19200, 19576, 23205, 24444, 25160, 24689, 23668, 23182, 22962, 22909, 
    23098, 23529, 24430, 25754, 26850, 23068, 25733, 26616, 26248, 25780, 
    25214, 24676,
  18299, 18645, 22733, 24181, 25096, 24624, 23666, 23192, 22946, 22953, 
    23077, 23539, 24453, 25640, 26541, 22550, 25746, 26620, 26287, 25875, 
    25305, 24758,
  17431, 17782, 22284, 24000, 25018, 24613, 23651, 23176, 22992, 22960, 
    23164, 23589, 24429, 25663, 26972, 22103, 25690, 26538, 26234, 25840, 
    25243, 24686,
  16897, 17231, 22165, 23952, 25047, 24639, 23647, 23193, 22935, 22915, 
    23133, 23528, 24407, 25541, 27018, 21914, 25661, 26482, 26111, 25692, 
    25124, 24566,
  16947, 17255, 22218, 24025, 25017, 24587, 23586, 23186, 22965, 22999, 
    23126, 23604, 24517, 25653, 26670, 21923, 25613, 26415, 26114, 25514, 
    24999, 24441,
  17706, 17941, 22566, 24212, 25081, 24553, 23553, 23176, 22971, 23012, 
    23153, 23584, 24559, 25668, 26776, 22137, 25596, 26499, 26088, 25622, 
    25045, 24489,
  19008, 19174, 23324, 24584, 25141, 24513, 23493, 23097, 22969, 22916, 
    23102, 23622, 24494, 25782, 27115, 22914, 25823, 26435, 26063, 25605, 
    25012, 24450,
  20486, 20605, 24185, 25074, 25284, 24522, 23518, 23170, 22992, 23026, 
    23111, 23650, 24641, 25863, 26719, 24001, 26237, 26455, 26091, 25567, 
    24975, 24337,
  21717, 21835, 24727, 25335, 25322, 24490, 23492, 23136, 23011, 23003, 
    23206, 23625, 24484, 26103, 26840, 24550, 26250, 26459, 26022, 25554, 
    25045, 24306,
  22487, 22599, 24884, 25358, 25237, 24411, 23479, 23123, 23004, 23051, 
    23097, 23557, 24501, 25991, 27054, 24520, 26238, 26517, 26151, 25635, 
    25058, 24514,
  22816, 22912, 24922, 25407, 25256, 24374, 23475, 23086, 23023, 22992, 
    23172, 23707, 24706, 26147, 26460, 24405, 26172, 26445, 26095, 25615, 
    25059, 24561,
  22915, 22990, 24911, 25365, 25259, 24370, 23434, 23103, 23047, 22999, 
    23238, 23786, 24721, 26038, 27026, 24335, 26225, 26438, 26060, 25590, 
    24977, 24461,
  22994, 23059, 25022, 25397, 25203, 24353, 23429, 23078, 22998, 23028, 
    23215, 23774, 24617, 25916, 27018, 24385, 26235, 26406, 25985, 25565, 
    25016, 24368,
  23138, 23216, 25123, 25426, 25182, 24273, 23375, 23106, 23004, 23022, 
    23240, 23700, 24650, 25971, 27301, 24574, 26379, 26324, 25876, 25498, 
    24820, 24335,
  23305, 23410, 25133, 25452, 25155, 24212, 23360, 23087, 22998, 22996, 
    23259, 23823, 24719, 26095, 27291, 24557, 26265, 26221, 25854, 25364, 
    24823, 24303,
  23422, 23550, 25193, 25488, 25097, 24211, 23335, 23104, 23050, 23116, 
    23354, 23843, 24784, 26087, 27291, 24390, 26185, 26201, 25768, 25337, 
    24749, 24192,
  23366, 23466, 25326, 25513, 25080, 24113, 23308, 23100, 23039, 23071, 
    23275, 23695, 24879, 26338, 27339, 24465, 26334, 26122, 25717, 25204, 
    24673, 24115,
  23077, 23057, 25462, 25567, 25022, 24054, 23277, 23115, 23054, 23055, 
    23266, 23847, 24872, 26066, 27109, 24465, 26285, 26141, 25663, 25237, 
    24645, 24125,
  22617, 22458, 25471, 25491, 24968, 24009, 23249, 23088, 23001, 23021, 
    23369, 23904, 25032, 26244, 27246, 24457, 26351, 26144, 25728, 25228, 
    24616, 24015,
  22399, 22160, 25480, 25459, 24878, 23924, 23227, 23050, 23014, 23077, 
    23301, 23918, 25033, 26484, 26960, 24394, 26403, 26119, 25756, 25204, 
    24591, 24017,
  27829, 27755, 27917, 27243, 25876, 24185, 22778, 22308, 22211, 22501, 
    23000, 23666, 24653, 25911, 26948, 28669, 28696, 27440, 26772, 25942, 
    24893, 23922,
  27829, 27767, 27883, 27207, 25954, 24249, 22833, 22314, 22231, 22540, 
    22927, 23637, 24641, 25822, 26732, 28531, 28505, 27207, 26400, 25700, 
    24676, 23842,
  27818, 27802, 27765, 27234, 26037, 24448, 22923, 22402, 22218, 22522, 
    23033, 23595, 24583, 25783, 26618, 28298, 28106, 26863, 26126, 25483, 
    24526, 23709,
  27747, 27793, 27694, 27249, 26072, 24501, 23010, 22432, 22259, 22506, 
    22931, 23583, 24639, 25831, 26779, 28149, 27839, 26552, 25847, 25228, 
    24487, 23689,
  27684, 27751, 27638, 27179, 26138, 24621, 23084, 22444, 22259, 22545, 
    22968, 23618, 24726, 25772, 26922, 27968, 27651, 26397, 25689, 25153, 
    24412, 23708,
  27591, 27630, 27500, 27122, 26119, 24637, 23104, 22562, 22261, 22546, 
    22947, 23603, 24586, 25876, 26694, 27861, 27451, 26328, 25697, 25228, 
    24481, 23880,
  27445, 27422, 27244, 26944, 26074, 24650, 23206, 22548, 22302, 22515, 
    22893, 23582, 24651, 25889, 26982, 27437, 27141, 26244, 25737, 25184, 
    24513, 23787,
  27235, 27175, 26932, 26672, 25957, 24646, 23228, 22610, 22305, 22529, 
    22918, 23546, 24502, 25524, 26675, 26833, 26641, 26026, 25679, 25222, 
    24463, 23860,
  27380, 27249, 26646, 26387, 25728, 24629, 23221, 22550, 22277, 22471, 
    22885, 23514, 24291, 25757, 26732, 26201, 25337, 25346, 25192, 24812, 
    24287, 23740,
  27128, 27005, 26404, 26231, 25746, 24635, 23293, 22585, 22210, 22474, 
    22879, 23499, 24416, 25437, 26660, 25641, 23485, 24480, 24771, 24650, 
    24217, 23706,
  26973, 26843, 26428, 26260, 25757, 24727, 23352, 22617, 22327, 22516, 
    22768, 23471, 24453, 25656, 26598, 25818, 24790, 25107, 25053, 24755, 
    24229, 23752,
  26949, 26825, 26595, 26385, 25834, 24783, 23377, 22623, 22314, 22556, 
    22830, 23551, 24359, 25493, 26865, 26278, 25809, 25540, 25287, 24867, 
    24312, 23618,
  26647, 26684, 26596, 26581, 26069, 24913, 23476, 22762, 22430, 22577, 
    22818, 23429, 24312, 25794, 26519, 26563, 26327, 25829, 25467, 25022, 
    24432, 23770,
  26791, 26879, 26779, 26712, 26204, 24972, 23563, 22785, 22426, 22524, 
    22949, 23477, 24461, 25697, 26525, 26928, 26753, 26041, 25546, 25100, 
    24398, 23875,
  26929, 27039, 26882, 26792, 26219, 25032, 23562, 22849, 22452, 22518, 
    22899, 23458, 24275, 25415, 26650, 27065, 26656, 25865, 25488, 24998, 
    24395, 23844,
  27020, 27113, 26888, 26822, 26224, 25061, 23619, 22866, 22484, 22560, 
    22938, 23431, 24419, 25632, 26669, 27097, 26613, 25857, 25437, 24933, 
    24381, 23801,
  27028, 27112, 26889, 26806, 26276, 25059, 23658, 22897, 22518, 22512, 
    22777, 23386, 24340, 25765, 26927, 27130, 26599, 25887, 25396, 24963, 
    24398, 23846,
  26969, 27061, 26809, 26729, 26263, 25104, 23637, 22920, 22509, 22604, 
    22868, 23479, 24384, 25641, 26896, 27079, 26462, 25799, 25340, 24894, 
    24396, 23864,
  26868, 26973, 26840, 26713, 26297, 25169, 23713, 22970, 22546, 22575, 
    22868, 23392, 24374, 25624, 26518, 27105, 26595, 25878, 25478, 24923, 
    24427, 23856,
  26753, 26846, 26741, 26721, 26296, 25176, 23734, 22970, 22534, 22539, 
    22992, 23455, 24119, 25482, 26563, 27169, 26874, 26167, 25684, 25183, 
    24496, 23930,
  26618, 26695, 26726, 26693, 26301, 25154, 23742, 23000, 22560, 22584, 
    22815, 23482, 24255, 25350, 26669, 27144, 26950, 26319, 25769, 25316, 
    24618, 23877,
  26467, 26543, 26672, 26626, 26214, 25178, 23783, 23038, 22608, 22600, 
    22812, 23345, 24281, 25419, 26626, 27076, 26741, 26266, 25816, 25316, 
    24693, 23943,
  26331, 26424, 26532, 26556, 26228, 25215, 23824, 23031, 22604, 22585, 
    22964, 23390, 24307, 25445, 26832, 27016, 26856, 26412, 25943, 25396, 
    24706, 24042,
  26261, 26382, 26538, 26612, 26282, 25248, 23844, 23036, 22595, 22590, 
    22940, 23401, 24349, 25472, 26568, 27088, 27119, 26523, 26013, 25357, 
    24737, 23994,
  26302, 26429, 26599, 26611, 26339, 25277, 23886, 23090, 22595, 22578, 
    22890, 23425, 24365, 25344, 26554, 27225, 27156, 26491, 25971, 25314, 
    24690, 24045,
  26440, 26554, 26644, 26684, 26329, 25317, 23901, 23094, 22643, 22600, 
    22887, 23401, 24205, 25367, 26987, 27210, 27184, 26525, 26068, 25467, 
    24790, 24076,
  26610, 26697, 26774, 26682, 26241, 25278, 23891, 23108, 22668, 22591, 
    22920, 23286, 24311, 25307, 26565, 27116, 27074, 26503, 26071, 25521, 
    24744, 24101,
  26728, 26789, 26744, 26673, 26240, 25287, 23963, 23133, 22693, 22585, 
    22835, 23322, 24304, 25582, 26718, 27107, 26924, 26524, 26144, 25643, 
    24857, 24095,
  26731, 26767, 26775, 26719, 26282, 25273, 23975, 23138, 22673, 22582, 
    22968, 23372, 24170, 25322, 26527, 27195, 27262, 26713, 26188, 25641, 
    24926, 24168,
  26599, 26620, 26751, 26697, 26300, 25326, 23960, 23126, 22675, 22564, 
    22865, 23315, 24374, 25456, 26405, 27254, 27396, 26775, 26351, 25784, 
    25015, 24335,
  26363, 26387, 26628, 26589, 26325, 25328, 23972, 23179, 22736, 22596, 
    22917, 23345, 24269, 25403, 26171, 27176, 27376, 26843, 26403, 25844, 
    25116, 24343,
  26094, 26135, 26532, 26513, 26218, 25293, 23973, 23196, 22692, 22610, 
    22898, 23375, 24339, 25287, 26604, 27053, 27320, 26825, 26381, 25925, 
    25194, 24443,
  25833, 25885, 26323, 26391, 26192, 25281, 24026, 23212, 22773, 22676, 
    22849, 23353, 24185, 25246, 26463, 26945, 27153, 26707, 26360, 25899, 
    25270, 24570,
  25577, 25628, 26235, 26320, 26132, 25273, 23998, 23215, 22749, 22674, 
    22906, 23375, 24179, 25475, 26650, 26828, 27066, 26749, 26351, 25919, 
    25321, 24604,
  25304, 25370, 26173, 26229, 26067, 25275, 23973, 23232, 22749, 22656, 
    22894, 23411, 24225, 25492, 26386, 26701, 26992, 26703, 26325, 25864, 
    25345, 24644,
  25034, 25136, 25924, 26124, 26004, 25262, 24019, 23253, 22774, 22625, 
    22824, 23351, 24137, 25503, 26487, 26582, 26944, 26629, 26262, 25857, 
    25313, 24656,
  24831, 24960, 25792, 26006, 25994, 25242, 23990, 23243, 22762, 22608, 
    22847, 23343, 24262, 25468, 26123, 26394, 26849, 26541, 26303, 25882, 
    25358, 24679,
  24745, 24849, 25547, 25925, 25949, 25180, 24000, 23235, 22799, 22665, 
    22785, 23399, 24100, 25401, 26819, 26196, 26635, 26440, 26088, 25758, 
    25179, 24692,
  24752, 24805, 25579, 25913, 25891, 25213, 23987, 23254, 22764, 22656, 
    22854, 23258, 24187, 25429, 26114, 26052, 26562, 26341, 25985, 25651, 
    25205, 24728,
  24778, 24796, 25761, 25998, 25938, 25227, 24066, 23269, 22770, 22674, 
    22847, 23390, 24133, 25479, 26249, 26035, 26606, 26365, 26034, 25713, 
    25250, 24656,
  24754, 24781, 25705, 26035, 25983, 25265, 24031, 23305, 22787, 22657, 
    22919, 23359, 24195, 25352, 26640, 25984, 26554, 26204, 25936, 25582, 
    25174, 24603,
  24695, 24758, 25615, 25990, 26005, 25254, 24021, 23271, 22836, 22671, 
    22923, 23429, 24171, 25311, 26288, 25817, 26650, 26363, 25991, 25644, 
    25131, 24638,
  24688, 24797, 25549, 25939, 26009, 25239, 24003, 23272, 22805, 22700, 
    22901, 23334, 24199, 25256, 26579, 25662, 26740, 26388, 26018, 25646, 
    25264, 24740,
  24820, 24953, 25649, 25999, 26049, 25297, 24048, 23273, 22864, 22646, 
    22888, 23287, 24306, 25330, 26362, 25750, 26741, 26407, 25993, 25565, 
    25106, 24699,
  25067, 25199, 25850, 26146, 26079, 25336, 24027, 23278, 22806, 22623, 
    22892, 23304, 24332, 25614, 26542, 25887, 26887, 26486, 26067, 25590, 
    25130, 24578,
  25325, 25440, 26022, 26270, 26161, 25284, 24037, 23297, 22822, 22684, 
    22913, 23264, 24251, 25389, 26521, 26020, 26862, 26435, 26029, 25573, 
    25074, 24504,
  25459, 25580, 26209, 26368, 26144, 25305, 23987, 23337, 22839, 22663, 
    22975, 23321, 24231, 25383, 26096, 26207, 26819, 26353, 25896, 25438, 
    24934, 24476,
  25436, 25597, 26181, 26351, 26162, 25259, 24037, 23304, 22837, 22689, 
    22940, 23342, 24128, 25235, 26254, 26222, 26690, 26304, 25809, 25407, 
    24862, 24407,
  25318, 25537, 26138, 26354, 26181, 25301, 24075, 23324, 22830, 22698, 
    22906, 23357, 24309, 25343, 26606, 26172, 26850, 26375, 25832, 25435, 
    24900, 24506,
  25222, 25458, 26057, 26279, 26099, 25348, 24029, 23325, 22880, 22732, 
    22992, 23337, 24155, 25276, 26531, 26031, 26916, 26516, 25976, 25526, 
    24830, 24319,
  25199, 25402, 25947, 26171, 26115, 25281, 24028, 23359, 22828, 22694, 
    23001, 23294, 24290, 25436, 26358, 25923, 26824, 26540, 26007, 25466, 
    24842, 24372,
  25231, 25381, 25937, 26230, 26101, 25310, 24059, 23336, 22876, 22754, 
    23000, 23357, 24085, 25321, 26485, 25883, 26724, 26529, 25901, 25407, 
    24816, 24293,
  25217, 25363, 26041, 26248, 26113, 25268, 24033, 23306, 22844, 22773, 
    22949, 23403, 24099, 25549, 26199, 26005, 26793, 26407, 25938, 25434, 
    24791, 24212,
  25064, 25258, 26066, 26251, 26082, 25262, 24007, 23352, 22892, 22782, 
    22990, 23362, 24129, 25271, 26197, 26086, 26963, 26451, 25900, 25430, 
    24817, 24151,
  24760, 25014, 25822, 26137, 26041, 25288, 24001, 23331, 22918, 22729, 
    22985, 23476, 24058, 25137, 26644, 25847, 26975, 26575, 26038, 25461, 
    24836, 24207,
  24334, 24618, 25633, 25978, 25961, 25253, 24010, 23320, 22874, 22701, 
    22935, 23408, 24327, 25305, 26816, 25494, 26744, 26688, 26234, 25592, 
    24855, 24233,
  23791, 24067, 25290, 25728, 25903, 25199, 24022, 23282, 22940, 22734, 
    22952, 23408, 24307, 25497, 26471, 25214, 26956, 26831, 26247, 25625, 
    24893, 24207,
  23069, 23329, 24876, 25505, 25804, 25203, 24006, 23332, 22893, 22771, 
    22953, 23411, 24241, 25425, 26614, 24921, 26834, 26863, 26288, 25713, 
    24912, 24281,
  22088, 22390, 24648, 25322, 25681, 25120, 24028, 23295, 22898, 22731, 
    22978, 23359, 24211, 25341, 26502, 24602, 26613, 26855, 26357, 25805, 
    25054, 24375,
  20872, 21273, 24424, 25221, 25634, 25134, 23953, 23283, 22900, 22769, 
    22892, 23397, 24306, 25563, 26525, 24421, 26540, 26946, 26453, 25838, 
    25176, 24415,
  19643, 20145, 23654, 24711, 25433, 25084, 23950, 23293, 22909, 22827, 
    22978, 23489, 24275, 25541, 26343, 23570, 26218, 26879, 26429, 25904, 
    25101, 24470,
  18713, 19279, 22593, 24024, 25126, 24970, 23968, 23293, 22917, 22786, 
    23015, 23420, 24177, 25503, 26546, 22177, 25101, 26601, 26404, 25875, 
    25154, 24451,
  18341, 18921, 22461, 23965, 25093, 24974, 23903, 23303, 22879, 22761, 
    23068, 23367, 24341, 25515, 26513, 22110, 25251, 26679, 26459, 26007, 
    25212, 24488,
  18589, 19124, 22758, 24148, 25121, 24945, 23903, 23292, 22906, 22815, 
    23068, 23519, 24278, 25551, 26862, 22581, 25493, 26713, 26446, 26026, 
    25270, 24557,
  19267, 19718, 23088, 24273, 25186, 24926, 23883, 23237, 22944, 22813, 
    23047, 23456, 24425, 25458, 26537, 22839, 25500, 26662, 26446, 26000, 
    25346, 24631,
  20069, 20422, 23537, 24600, 25313, 24939, 23897, 23260, 22939, 22856, 
    23070, 23399, 24252, 25408, 27038, 23386, 25654, 26726, 26456, 26044, 
    25321, 24651,
  20743, 21031, 23965, 24836, 25378, 24917, 23843, 23252, 22980, 22818, 
    22981, 23458, 24366, 25374, 26558, 23863, 25932, 26689, 26459, 26006, 
    25298, 24644,
  21181, 21467, 24009, 24829, 25381, 24888, 23826, 23247, 22899, 22768, 
    23112, 23483, 24251, 25454, 26592, 23887, 25944, 26714, 26425, 25983, 
    25253, 24714,
  21421, 21733, 23935, 24774, 25349, 24872, 23829, 23237, 22906, 22840, 
    22984, 23463, 24200, 25489, 26815, 23761, 25793, 26659, 26334, 25899, 
    25267, 24682,
  21552, 21851, 23949, 24826, 25303, 24902, 23828, 23279, 22905, 22847, 
    23124, 23426, 24362, 25581, 26744, 23788, 25804, 26625, 26332, 25791, 
    25128, 24489,
  21611, 21860, 24152, 24936, 25351, 24870, 23760, 23221, 22924, 22834, 
    23021, 23432, 24320, 25370, 26697, 23874, 25770, 26601, 26235, 25824, 
    25176, 24544,
  21600, 21812, 24193, 25022, 25368, 24833, 23751, 23232, 22972, 22826, 
    23042, 23466, 24320, 25479, 26526, 24038, 25762, 26599, 26313, 25753, 
    25106, 24494,
  21502, 21738, 24114, 24992, 25347, 24796, 23749, 23242, 22950, 22949, 
    23054, 23478, 24380, 25452, 26683, 24075, 25965, 26612, 26236, 25723, 
    25165, 24656,
  21311, 21605, 24047, 24936, 25346, 24783, 23759, 23235, 22962, 22907, 
    23036, 23498, 24418, 25740, 26699, 24115, 26094, 26587, 26186, 25788, 
    25141, 24617,
  20991, 21348, 23978, 24876, 25336, 24727, 23693, 23193, 22949, 22893, 
    23085, 23468, 24321, 25787, 26663, 24024, 26117, 26628, 26228, 25816, 
    25187, 24598,
  20514, 20888, 23824, 24845, 25268, 24744, 23682, 23193, 22956, 22949, 
    23166, 23472, 24461, 25537, 26834, 23842, 25930, 26590, 26269, 25818, 
    25296, 24727,
  19837, 20213, 23584, 24684, 25203, 24659, 23685, 23189, 23004, 22841, 
    23125, 23519, 24536, 25750, 26871, 23507, 25888, 26581, 26263, 25863, 
    25292, 24853,
  19006, 19373, 23033, 24389, 25150, 24653, 23670, 23214, 22956, 23029, 
    23112, 23511, 24424, 25806, 26826, 22967, 25788, 26491, 26233, 25797, 
    25242, 24774,
  18160, 18535, 22511, 24159, 25076, 24643, 23621, 23162, 22945, 22958, 
    23036, 23533, 24534, 25685, 26799, 22260, 25565, 26524, 26200, 25743, 
    25219, 24741,
  17594, 17936, 22225, 24017, 24992, 24576, 23629, 23185, 22953, 22931, 
    23089, 23607, 24512, 25742, 26867, 21913, 25506, 26476, 26147, 25788, 
    25176, 24583,
  17566, 17852, 22326, 24095, 25001, 24627, 23637, 23179, 22966, 22922, 
    23070, 23609, 24443, 25807, 26521, 21868, 25452, 26460, 26095, 25666, 
    24962, 24350,
  18202, 18393, 22530, 24226, 25011, 24558, 23606, 23154, 22980, 23001, 
    23134, 23645, 24571, 25729, 26659, 22005, 25571, 26506, 26138, 25631, 
    24995, 24445,
  19350, 19462, 23183, 24539, 25149, 24494, 23545, 23146, 23020, 23010, 
    23214, 23690, 24553, 25712, 26796, 22732, 25722, 26472, 26091, 25664, 
    25097, 24473,
  20673, 20740, 24096, 25001, 25229, 24520, 23592, 23154, 22996, 23004, 
    23175, 23683, 24480, 25897, 26734, 23771, 26063, 26464, 26153, 25725, 
    25129, 24540,
  21787, 21860, 24714, 25287, 25335, 24458, 23534, 23134, 23026, 23004, 
    23162, 23686, 24601, 25682, 26729, 24418, 26237, 26461, 26196, 25744, 
    25204, 24663,
  22502, 22575, 24870, 25383, 25290, 24463, 23503, 23135, 22978, 23000, 
    23183, 23715, 24427, 26025, 26828, 24529, 26282, 26475, 26125, 25806, 
    25237, 24651,
  22827, 22891, 24868, 25399, 25335, 24425, 23462, 23134, 23030, 23014, 
    23121, 23723, 24459, 25950, 27069, 24455, 26191, 26468, 26123, 25730, 
    25232, 24751,
  22938, 22993, 25009, 25422, 25243, 24377, 23452, 23113, 23019, 23012, 
    23224, 23606, 24642, 25741, 26950, 24415, 26268, 26432, 26164, 25723, 
    25290, 24651,
  23020, 23075, 25014, 25446, 25230, 24284, 23418, 23143, 23034, 23032, 
    23157, 23711, 24698, 26145, 27057, 24449, 26315, 26421, 26022, 25635, 
    25144, 24591,
  23162, 23224, 25076, 25475, 25201, 24274, 23431, 23128, 23054, 23046, 
    23220, 23804, 24864, 26019, 27001, 24478, 26316, 26325, 26001, 25631, 
    25012, 24478,
  23347, 23414, 25153, 25552, 25165, 24200, 23399, 23129, 23060, 23089, 
    23288, 23803, 24655, 26258, 26956, 24516, 26282, 26280, 25889, 25591, 
    24983, 24420,
  23514, 23589, 25329, 25512, 25115, 24184, 23335, 23105, 23033, 23031, 
    23235, 23780, 24762, 25887, 27185, 24459, 26278, 26246, 25837, 25396, 
    24768, 24322,
  23534, 23589, 25400, 25562, 25084, 24114, 23281, 23107, 23060, 23030, 
    23415, 23839, 24765, 26067, 27021, 24636, 26282, 26189, 25717, 25250, 
    24707, 24212,
  23325, 23287, 25510, 25598, 25058, 24079, 23291, 23143, 23067, 23028, 
    23321, 23837, 24813, 26129, 27171, 24690, 26341, 26100, 25657, 25197, 
    24672, 24175,
  22925, 22776, 25520, 25540, 24967, 23974, 23242, 23115, 23070, 23071, 
    23293, 23953, 24891, 26166, 27121, 24662, 26313, 26044, 25612, 25224, 
    24649, 24018,
  22729, 22510, 25582, 25549, 24893, 23911, 23203, 23084, 23047, 23050, 
    23356, 23909, 24971, 26165, 27312, 24572, 26291, 26071, 25632, 25182, 
    24548, 24040,
  27748, 27628, 27878, 27188, 25857, 24167, 22780, 22328, 22185, 22518, 
    23094, 23654, 24732, 25755, 26769, 28568, 28326, 27045, 26384, 25618, 
    24583, 23721,
  27738, 27628, 27794, 27176, 25935, 24272, 22842, 22351, 22237, 22605, 
    22979, 23546, 24629, 25701, 26674, 28369, 28086, 26739, 26123, 25407, 
    24545, 23760,
  27709, 27639, 27666, 27116, 25979, 24361, 22967, 22406, 22270, 22585, 
    22979, 23615, 24682, 26064, 26762, 28132, 27735, 26497, 25863, 25240, 
    24401, 23634,
  27628, 27621, 27556, 27103, 26022, 24468, 23009, 22446, 22300, 22502, 
    22986, 23599, 24404, 25707, 26995, 27932, 27488, 26236, 25584, 24965, 
    24337, 23600,
  27569, 27590, 27507, 27066, 26085, 24545, 23094, 22508, 22265, 22568, 
    23014, 23604, 24367, 25788, 26603, 27814, 27488, 26291, 25660, 25051, 
    24350, 23592,
  27487, 27491, 27432, 27011, 26082, 24564, 23103, 22508, 22288, 22512, 
    22901, 23543, 24456, 25690, 26862, 27657, 27423, 26344, 25799, 25109, 
    24393, 23712,
  27354, 27308, 27132, 26828, 25984, 24617, 23215, 22532, 22334, 22514, 
    22851, 23544, 24467, 25657, 26901, 27242, 27057, 26210, 25735, 25133, 
    24452, 23759,
  27163, 27094, 26820, 26534, 25910, 24648, 23195, 22560, 22308, 22538, 
    22890, 23648, 24537, 25459, 26448, 26487, 26415, 25978, 25568, 25139, 
    24502, 23878,
  27333, 27212, 26562, 26346, 25690, 24587, 23244, 22572, 22245, 22516, 
    22800, 23489, 24472, 25579, 27014, 25957, 24762, 25138, 25129, 24786, 
    24257, 23812,
  27104, 27015, 26485, 26260, 25698, 24676, 23310, 22611, 22257, 22476, 
    22939, 23520, 24543, 25533, 26519, 25824, 23911, 24763, 24901, 24773, 
    24314, 23745,
  26959, 26877, 26531, 26338, 25787, 24730, 23368, 22584, 22274, 22524, 
    22882, 23506, 24572, 25493, 26285, 26156, 25166, 25282, 25114, 24884, 
    24289, 23791,
  26933, 26846, 26647, 26443, 25870, 24760, 23393, 22648, 22323, 22432, 
    22867, 23390, 24382, 25523, 26167, 26541, 25595, 25461, 25238, 24859, 
    24313, 23777,
  26617, 26663, 26638, 26584, 26079, 24933, 23493, 22767, 22433, 22547, 
    22898, 23515, 24473, 25599, 26590, 26638, 26200, 25751, 25424, 25033, 
    24390, 23889,
  26744, 26821, 26765, 26650, 26171, 24955, 23520, 22793, 22446, 22521, 
    22898, 23552, 24539, 25580, 26857, 26931, 26837, 26070, 25572, 25049, 
    24508, 23940,
  26879, 26970, 26884, 26765, 26187, 25057, 23567, 22837, 22476, 22572, 
    22877, 23482, 24340, 25619, 26784, 27094, 26997, 26250, 25679, 25133, 
    24492, 23876,
  26987, 27056, 26895, 26781, 26208, 25033, 23625, 22871, 22460, 22557, 
    22875, 23477, 24326, 25500, 26447, 27128, 26747, 25937, 25539, 24969, 
    24370, 23847,
  27024, 27077, 26913, 26760, 26253, 25118, 23667, 22908, 22540, 22557, 
    22871, 23392, 24320, 25515, 26574, 27100, 26367, 25657, 25298, 24868, 
    24348, 23804,
  26984, 27045, 26816, 26753, 26254, 25040, 23675, 22911, 22546, 22526, 
    22905, 23502, 24326, 25424, 26506, 27047, 26441, 25678, 25325, 24936, 
    24392, 23870,
  26872, 26963, 26775, 26772, 26256, 25149, 23715, 22951, 22526, 22557, 
    22879, 23479, 24365, 25435, 26436, 27072, 26699, 25929, 25477, 25065, 
    24390, 23848,
  26718, 26819, 26755, 26699, 26229, 25153, 23705, 22948, 22548, 22543, 
    22896, 23387, 24357, 25559, 26544, 27134, 26990, 26204, 25663, 25213, 
    24556, 23949,
  26529, 26625, 26713, 26641, 26217, 25168, 23754, 22990, 22592, 22555, 
    22838, 23396, 24354, 25485, 26547, 27103, 26917, 26341, 25850, 25383, 
    24632, 24043,
  26331, 26417, 26578, 26522, 26181, 25119, 23806, 23011, 22637, 22559, 
    22821, 23553, 24363, 25763, 26656, 26918, 26607, 26260, 25878, 25383, 
    24682, 24109,
  26164, 26252, 26526, 26515, 26187, 25207, 23806, 23026, 22662, 22582, 
    22842, 23378, 24345, 25601, 26559, 26813, 26429, 26247, 25907, 25426, 
    24696, 23974,
  26077, 26182, 26426, 26511, 26212, 25268, 23887, 23085, 22650, 22554, 
    22867, 23488, 24346, 25412, 26584, 26915, 26768, 26394, 25971, 25399, 
    24720, 24026,
  26106, 26211, 26545, 26601, 26278, 25252, 23878, 23068, 22662, 22626, 
    22884, 23408, 24297, 25370, 26674, 27095, 27085, 26579, 26051, 25542, 
    24793, 24097,
  26230, 26316, 26631, 26624, 26239, 25262, 23893, 23111, 22662, 22596, 
    22984, 23485, 24208, 25320, 26397, 27066, 27051, 26547, 26065, 25626, 
    24856, 24176,
  26384, 26439, 26633, 26588, 26235, 25259, 23907, 23157, 22650, 22570, 
    22895, 23367, 24211, 25462, 26695, 27012, 26922, 26562, 26187, 25618, 
    24873, 24187,
  26493, 26527, 26616, 26613, 26270, 25251, 23889, 23140, 22679, 22602, 
    22935, 23409, 24231, 25419, 26615, 26985, 26935, 26568, 26128, 25666, 
    24961, 24226,
  26507, 26524, 26678, 26637, 26276, 25262, 23936, 23140, 22637, 22642, 
    22922, 23403, 24348, 25264, 26564, 27057, 27228, 26693, 26201, 25682, 
    25036, 24307,
  26418, 26421, 26688, 26635, 26322, 25341, 23942, 23149, 22701, 22650, 
    22836, 23320, 24243, 25414, 26615, 27082, 27300, 26725, 26301, 25788, 
    25087, 24481,
  26261, 26256, 26447, 26550, 26203, 25266, 23964, 23196, 22733, 22578, 
    22886, 23437, 24247, 25356, 26613, 27046, 27342, 26822, 26375, 25966, 
    25202, 24570,
  26098, 26094, 26365, 26456, 26229, 25274, 23979, 23180, 22733, 22626, 
    22876, 23315, 24125, 25336, 26372, 26898, 27304, 26762, 26393, 25966, 
    25253, 24550,
  25945, 25953, 26335, 26443, 26176, 25296, 23970, 23211, 22734, 22638, 
    22832, 23455, 24261, 25421, 26338, 26817, 27213, 26781, 26338, 25909, 
    25310, 24570,
  25777, 25801, 26296, 26349, 26149, 25281, 23959, 23240, 22760, 22597, 
    22872, 23337, 24226, 25291, 26647, 26706, 27013, 26707, 26301, 25899, 
    25304, 24630,
  25566, 25620, 26063, 26269, 26097, 25263, 23989, 23240, 22775, 22598, 
    23006, 23421, 24314, 25336, 26440, 26610, 27051, 26675, 26260, 25912, 
    25303, 24698,
  25331, 25421, 25957, 26177, 26082, 25293, 23980, 23261, 22754, 22697, 
    22915, 23339, 24340, 25510, 26329, 26452, 26916, 26573, 26191, 25900, 
    25334, 24763,
  25140, 25248, 25766, 26062, 26010, 25264, 23999, 23280, 22846, 22654, 
    22915, 23397, 24329, 25357, 26675, 26222, 26903, 26528, 26178, 25837, 
    25410, 24739,
  25046, 25129, 25543, 25922, 25924, 25220, 23979, 23281, 22793, 22673, 
    22862, 23448, 24207, 25471, 26825, 25938, 26771, 26419, 26066, 25787, 
    25321, 24746,
  25038, 25086, 25641, 25945, 25938, 25230, 24021, 23288, 22811, 22692, 
    22814, 23368, 24287, 25266, 26870, 25855, 26591, 26371, 26081, 25798, 
    25385, 24781,
  25062, 25096, 25750, 26081, 25974, 25233, 24016, 23254, 22799, 22646, 
    22915, 23345, 24129, 25236, 26176, 25947, 26559, 26359, 25985, 25674, 
    25322, 24796,
  25063, 25119, 25805, 26099, 26001, 25223, 23956, 23260, 22776, 22619, 
    22916, 23407, 24142, 25268, 26484, 25959, 26671, 26365, 25997, 25699, 
    25336, 24951,
  25054, 25143, 25672, 26032, 26034, 25254, 24011, 23258, 22827, 22660, 
    22886, 23392, 24158, 25307, 26632, 25801, 26816, 26466, 26045, 25754, 
    25413, 24953,
  25105, 25232, 25424, 25957, 25973, 25303, 24006, 23333, 22807, 22643, 
    22964, 23367, 24197, 25307, 26375, 25526, 26632, 26462, 26086, 25743, 
    25324, 24879,
  25278, 25423, 25633, 26081, 26068, 25345, 24001, 23272, 22823, 22674, 
    22880, 23298, 24126, 25588, 26557, 25606, 26659, 26444, 25985, 25675, 
    25223, 24806,
  25521, 25670, 26031, 26283, 26161, 25338, 24054, 23277, 22853, 22769, 
    22807, 23376, 24244, 25378, 26484, 26018, 26940, 26516, 26045, 25638, 
    25286, 24778,
  25725, 25868, 26407, 26485, 26248, 25309, 23959, 23285, 22836, 22718, 
    22885, 23299, 24190, 25417, 26570, 26429, 27003, 26472, 25918, 25546, 
    25146, 24618,
  25781, 25936, 26429, 26481, 26204, 25319, 24027, 23325, 22848, 22696, 
    22926, 23335, 24239, 25381, 26333, 26537, 26872, 26347, 25847, 25449, 
    25018, 24495,
  25702, 25887, 26275, 26431, 26195, 25299, 24008, 23280, 22860, 22703, 
    22972, 23370, 24229, 25086, 26421, 26393, 26906, 26428, 25849, 25400, 
    24838, 24487,
  25573, 25800, 26200, 26324, 26165, 25301, 24021, 23299, 22827, 22749, 
    22947, 23446, 24221, 25336, 26787, 26295, 26946, 26426, 25929, 25403, 
    24806, 24339,
  25506, 25745, 26171, 26344, 26183, 25314, 24024, 23336, 22859, 22723, 
    22954, 23370, 24215, 25515, 26445, 26316, 26919, 26431, 25858, 25264, 
    24813, 24258,
  25528, 25746, 26218, 26369, 26179, 25340, 24010, 23293, 22856, 22708, 
    22954, 23350, 24193, 25441, 26556, 26325, 26878, 26353, 25861, 25340, 
    24780, 24318,
  25601, 25791, 26223, 26401, 26211, 25326, 24029, 23338, 22882, 22728, 
    22946, 23289, 24110, 25443, 26513, 26341, 26857, 26356, 25844, 25281, 
    24716, 24272,
  25619, 25830, 26240, 26368, 26126, 25291, 23997, 23302, 22837, 22627, 
    22890, 23325, 24283, 25474, 26466, 26380, 26989, 26459, 25964, 25326, 
    24755, 24272,
  25500, 25763, 26215, 26334, 26099, 25287, 24010, 23318, 22854, 22764, 
    22928, 23426, 24194, 25239, 26682, 26368, 27091, 26612, 26071, 25503, 
    24864, 24285,
  25221, 25522, 26100, 26279, 26091, 25246, 23990, 23303, 22859, 22717, 
    22973, 23383, 24232, 25351, 26419, 26291, 27153, 26676, 26168, 25528, 
    24825, 24226,
  24781, 25078, 25922, 26115, 26034, 25228, 24016, 23354, 22901, 22735, 
    23009, 23419, 24308, 25315, 26519, 26069, 27153, 26782, 26260, 25653, 
    24895, 24259,
  24162, 24434, 25579, 25925, 25959, 25258, 23962, 23299, 22882, 22765, 
    23046, 23431, 24193, 25378, 26612, 25690, 27034, 26825, 26238, 25692, 
    25010, 24319,
  23331, 23591, 25031, 25601, 25850, 25242, 24001, 23293, 22921, 22734, 
    22959, 23446, 24210, 25474, 26596, 25046, 26658, 26829, 26328, 25766, 
    25048, 24394,
  22270, 22588, 24593, 25364, 25706, 25163, 23982, 23303, 22901, 22757, 
    22942, 23423, 24360, 25401, 26364, 24472, 26331, 26856, 26453, 25946, 
    25139, 24528,
  21063, 21481, 24217, 25147, 25656, 25084, 23948, 23294, 22928, 22795, 
    23035, 23410, 24302, 25374, 26485, 24341, 26574, 26925, 26472, 25954, 
    25229, 24635,
  19939, 20446, 23540, 24715, 25395, 25072, 23939, 23286, 22876, 22815, 
    23035, 23431, 24118, 25543, 27091, 23557, 26141, 26807, 26422, 25990, 
    25167, 24529,
  19171, 19724, 22740, 24107, 25147, 24987, 23932, 23287, 22902, 22763, 
    23073, 23560, 24325, 25445, 26537, 22386, 25160, 26631, 26332, 25979, 
    25270, 24577,
  18957, 19506, 22776, 24166, 25141, 24948, 23876, 23293, 22938, 22801, 
    22959, 23354, 24322, 25415, 26297, 22511, 25479, 26701, 26397, 25980, 
    25227, 24588,
  19295, 19788, 23142, 24389, 25206, 24920, 23887, 23301, 22926, 22832, 
    23036, 23459, 24404, 25455, 26378, 22968, 25715, 26707, 26458, 25968, 
    25292, 24676,
  19965, 20373, 23531, 24536, 25268, 24942, 23917, 23304, 22961, 22822, 
    23076, 23540, 24366, 25316, 26827, 23236, 25601, 26691, 26431, 26054, 
    25356, 24724,
  20667, 20994, 23949, 24804, 25378, 24944, 23854, 23246, 22907, 22838, 
    23008, 23437, 24309, 25480, 26568, 23804, 25963, 26749, 26565, 26048, 
    25407, 24790,
  21201, 21485, 24076, 24902, 25414, 24945, 23879, 23230, 22932, 22823, 
    23078, 23431, 24407, 25562, 26537, 24070, 26074, 26727, 26500, 26059, 
    25287, 24744,
  21515, 21805, 24010, 24939, 25351, 24941, 23846, 23231, 22922, 22864, 
    23155, 23516, 24364, 25750, 26936, 23977, 25949, 26701, 26418, 26000, 
    25281, 24700,
  21674, 21976, 23939, 24868, 25365, 24880, 23829, 23236, 22955, 22884, 
    23013, 23527, 24284, 25532, 26876, 23846, 25865, 26688, 26381, 25861, 
    25237, 24675,
  21751, 22021, 23991, 24895, 25381, 24874, 23776, 23243, 22963, 22861, 
    23041, 23498, 24420, 25412, 26557, 23847, 25783, 26584, 26254, 25814, 
    25207, 24609,
  21756, 21976, 24222, 25046, 25376, 24867, 23787, 23250, 22947, 22954, 
    23075, 23595, 24198, 25588, 26531, 24115, 25948, 26624, 26359, 25816, 
    25261, 24710,
  21685, 21888, 24301, 25081, 25423, 24853, 23781, 23243, 22972, 22853, 
    23076, 23508, 24297, 25588, 26743, 24348, 26127, 26650, 26326, 25807, 
    25306, 24741,
  21548, 21795, 24205, 25037, 25383, 24809, 23723, 23221, 22929, 22906, 
    23176, 23580, 24351, 25531, 26696, 24337, 26324, 26671, 26331, 25864, 
    25308, 24783,
  21377, 21686, 23970, 24914, 25310, 24802, 23769, 23205, 22971, 22893, 
    23167, 23481, 24337, 25675, 27110, 24168, 26185, 26638, 26316, 25906, 
    25386, 24817,
  21161, 21524, 23995, 24903, 25317, 24760, 23709, 23204, 22965, 22925, 
    23059, 23555, 24319, 25603, 26659, 24078, 26170, 26628, 26247, 25865, 
    25312, 24758,
  20858, 21239, 24041, 24921, 25278, 24713, 23698, 23176, 22953, 22940, 
    23092, 23512, 24438, 25719, 26979, 24099, 26176, 26620, 26261, 25897, 
    25286, 24800,
  20379, 20783, 23968, 24896, 25307, 24715, 23671, 23212, 22993, 22915, 
    23154, 23529, 24541, 25733, 26682, 23949, 26134, 26516, 26234, 25768, 
    25243, 24625,
  19727, 20144, 23570, 24701, 25200, 24737, 23672, 23257, 22964, 22931, 
    23218, 23537, 24580, 25689, 26579, 23458, 26022, 26565, 26190, 25807, 
    25232, 24740,
  19007, 19430, 22933, 24387, 25150, 24670, 23679, 23183, 23024, 22955, 
    23151, 23617, 24333, 25631, 26759, 22737, 25687, 26540, 26261, 25828, 
    25323, 24728,
  18490, 18851, 22675, 24253, 25105, 24631, 23621, 23167, 23009, 22956, 
    23163, 23666, 24414, 25539, 26475, 22245, 25534, 26426, 26152, 25774, 
    25101, 24529,
  18412, 18686, 22709, 24296, 25051, 24602, 23578, 23201, 22996, 22919, 
    23162, 23592, 24357, 25794, 26839, 22146, 25530, 26418, 26093, 25651, 
    25104, 24476,
  18900, 19064, 22800, 24347, 25101, 24541, 23591, 23173, 22960, 22978, 
    23128, 23630, 24529, 25659, 26491, 22106, 25407, 26443, 26095, 25574, 
    25048, 24451,
  19834, 19920, 23314, 24626, 25119, 24509, 23582, 23183, 23002, 23006, 
    23197, 23597, 24527, 25837, 26532, 22562, 25496, 26538, 26124, 25711, 
    25112, 24546,
  20932, 20984, 24042, 24979, 25187, 24472, 23521, 23183, 23016, 23000, 
    23197, 23740, 24659, 25951, 26766, 23485, 25824, 26443, 26152, 25767, 
    25187, 24601,
  21876, 21942, 24634, 25279, 25305, 24517, 23491, 23157, 22991, 23018, 
    23147, 23636, 24601, 25724, 26734, 24265, 26222, 26498, 26181, 25841, 
    25271, 24629,
  22505, 22579, 24824, 25379, 25295, 24468, 23492, 23170, 23025, 23026, 
    23183, 23637, 24635, 25651, 27104, 24465, 26329, 26462, 26117, 25823, 
    25304, 24717,
  22817, 22893, 24940, 25420, 25245, 24428, 23495, 23169, 23035, 23039, 
    23281, 23763, 24655, 26035, 27026, 24419, 26275, 26470, 26136, 25747, 
    25221, 24711,
  22950, 23029, 24995, 25449, 25259, 24390, 23462, 23159, 23042, 23062, 
    23264, 23796, 24751, 25776, 27149, 24407, 26321, 26412, 26107, 25672, 
    25114, 24577,
  23057, 23135, 25028, 25478, 25246, 24337, 23428, 23140, 23025, 23062, 
    23330, 23752, 24872, 25898, 27322, 24402, 26331, 26314, 25991, 25666, 
    25082, 24491,
  23219, 23282, 25179, 25480, 25196, 24290, 23423, 23169, 23033, 23074, 
    23235, 23751, 24823, 25834, 27250, 24493, 26240, 26291, 25953, 25543, 
    24944, 24397,
  23431, 23464, 25266, 25513, 25189, 24247, 23370, 23153, 23080, 23083, 
    23263, 23839, 24729, 26288, 27034, 24539, 26318, 26274, 25929, 25521, 
    24966, 24385,
  23637, 23658, 25354, 25538, 25132, 24179, 23341, 23161, 23080, 23059, 
    23301, 23824, 24859, 25996, 27249, 24533, 26312, 26262, 25871, 25487, 
    24846, 24267,
  23704, 23718, 25528, 25577, 25080, 24144, 23332, 23168, 23051, 23055, 
    23276, 23886, 24808, 26315, 27076, 24701, 26374, 26183, 25778, 25335, 
    24709, 24264,
  23536, 23498, 25529, 25588, 25025, 24064, 23332, 23125, 23087, 23073, 
    23293, 23812, 25060, 26212, 26993, 24801, 26369, 26094, 25662, 25184, 
    24629, 24114,
  23167, 23057, 25572, 25575, 24977, 24001, 23259, 23114, 23131, 23165, 
    23361, 23814, 24998, 26454, 27231, 24841, 26398, 26096, 25604, 25167, 
    24651, 24097,
  22982, 22819, 25516, 25531, 24943, 23939, 23288, 23080, 23079, 23121, 
    23382, 23851, 24954, 26100, 27362, 24757, 26357, 26007, 25542, 25020, 
    24499, 23958,
  27651, 27523, 27738, 27109, 25836, 24196, 22806, 22368, 22217, 22563, 
    22987, 23649, 24695, 25996, 26632, 28357, 27919, 26776, 26100, 25385, 
    24409, 23679,
  27632, 27507, 27653, 27034, 25881, 24261, 22875, 22338, 22255, 22511, 
    22958, 23635, 24666, 25847, 26696, 28063, 27684, 26557, 25921, 25242, 
    24504, 23733,
  27585, 27489, 27487, 27001, 25882, 24350, 22940, 22408, 22215, 22490, 
    22946, 23610, 24788, 25812, 26835, 27853, 27376, 26293, 25791, 25237, 
    24506, 23760,
  27494, 27456, 27395, 26951, 25921, 24399, 22957, 22453, 22245, 22534, 
    22965, 23569, 24528, 25728, 26557, 27712, 27279, 26205, 25671, 25104, 
    24385, 23793,
  27439, 27438, 27316, 26998, 25987, 24489, 23025, 22457, 22277, 22551, 
    22868, 23553, 24509, 25693, 26553, 27567, 27228, 26325, 25788, 25278, 
    24474, 23771,
  27371, 27371, 27210, 26943, 25990, 24579, 23121, 22487, 22285, 22560, 
    22916, 23632, 24567, 25773, 26446, 27423, 27357, 26392, 25866, 25192, 
    24518, 23905,
  27263, 27224, 26979, 26778, 25976, 24617, 23168, 22537, 22317, 22540, 
    22921, 23617, 24598, 25768, 26578, 26975, 27054, 26345, 25850, 25292, 
    24646, 24032,
  27527, 27386, 26723, 26421, 25743, 24540, 23190, 22498, 22251, 22522, 
    22841, 23497, 24447, 25489, 26879, 26429, 25828, 25648, 25450, 25050, 
    24503, 23885,
  27336, 27212, 26548, 26335, 25669, 24644, 23217, 22539, 22245, 22525, 
    22872, 23502, 24402, 25551, 26685, 25919, 24478, 24948, 25050, 24795, 
    24356, 23751,
  27143, 27059, 26563, 26345, 25731, 24646, 23314, 22574, 22286, 22493, 
    22866, 23456, 24242, 25657, 26510, 26220, 25492, 25424, 25264, 24931, 
    24381, 23837,
  26606, 26646, 26565, 26485, 25907, 24778, 23426, 22734, 22427, 22588, 
    22937, 23490, 24407, 25476, 26869, 26449, 26188, 25694, 25386, 24980, 
    24435, 23784,
  26560, 26604, 26581, 26529, 26019, 24817, 23440, 22779, 22436, 22505, 
    22896, 23429, 24374, 25666, 26764, 26522, 25799, 25553, 25267, 24933, 
    24376, 23856,
  26593, 26651, 26599, 26516, 26032, 24888, 23462, 22784, 22436, 22545, 
    22936, 23475, 24441, 25750, 26594, 26676, 26227, 25791, 25443, 24955, 
    24304, 23808,
  26690, 26761, 26673, 26655, 26182, 24986, 23528, 22818, 22449, 22560, 
    22953, 23592, 24489, 25589, 26874, 26949, 26709, 26011, 25570, 25064, 
    24397, 23892,
  26815, 26891, 26842, 26759, 26174, 25001, 23586, 22829, 22464, 22606, 
    22875, 23440, 24565, 25506, 27044, 27131, 26906, 26031, 25491, 25006, 
    24356, 23781,
  26934, 26985, 26856, 26759, 26193, 25025, 23598, 22867, 22446, 22560, 
    22931, 23434, 24213, 25768, 26967, 27121, 26481, 25618, 25254, 24779, 
    24233, 23758,
  26993, 27022, 26838, 26732, 26231, 25071, 23654, 22901, 22506, 22565, 
    22835, 23430, 24376, 25564, 26444, 27028, 26368, 25641, 25296, 24983, 
    24378, 23890,
  26967, 27000, 26791, 26647, 26222, 25100, 23714, 22918, 22543, 22583, 
    22855, 23382, 24389, 25533, 26613, 27050, 26705, 25963, 25468, 25051, 
    24376, 23728,
  26850, 26917, 26759, 26653, 26203, 25136, 23709, 22933, 22537, 22566, 
    22829, 23392, 24409, 25530, 26471, 27056, 26943, 26251, 25735, 25179, 
    24464, 23921,
  26669, 26754, 26720, 26612, 26145, 25104, 23706, 22971, 22578, 22587, 
    22932, 23428, 24277, 25596, 26747, 27065, 26968, 26332, 25784, 25272, 
    24535, 23841,
  26443, 26527, 26714, 26594, 26170, 25121, 23762, 23022, 22569, 22586, 
    22887, 23416, 24312, 25415, 26538, 26956, 26937, 26318, 25834, 25305, 
    24546, 23854,
  26210, 26284, 26466, 26544, 26155, 25193, 23803, 23051, 22629, 22585, 
    22860, 23444, 24402, 25270, 26456, 26793, 26616, 26229, 25785, 25262, 
    24610, 23861,
  26020, 26095, 26482, 26498, 26180, 25196, 23796, 23050, 22612, 22570, 
    22882, 23441, 24335, 25512, 26698, 26764, 26407, 26137, 25780, 25385, 
    24699, 23965,
  25920, 26012, 26429, 26481, 26214, 25204, 23826, 23090, 22656, 22572, 
    22954, 23417, 24387, 25511, 26550, 26907, 26869, 26414, 25975, 25396, 
    24723, 24019,
  25932, 26021, 26460, 26488, 26200, 25190, 23872, 23129, 22636, 22571, 
    22828, 23494, 24217, 25223, 26692, 27029, 27112, 26541, 26071, 25520, 
    24778, 24110,
  26024, 26087, 26528, 26524, 26215, 25160, 23890, 23125, 22665, 22619, 
    22915, 23480, 24272, 25376, 26663, 27004, 26996, 26503, 26104, 25524, 
    24929, 24154,
  26138, 26161, 26475, 26557, 26176, 25231, 23849, 23088, 22626, 22579, 
    22790, 23413, 24307, 25483, 26683, 26912, 26943, 26524, 26156, 25653, 
    24953, 24226,
  26213, 26214, 26435, 26485, 26166, 25235, 23908, 23123, 22697, 22668, 
    22848, 23330, 24181, 25410, 26691, 26897, 27024, 26552, 26106, 25626, 
    24946, 24200,
  26222, 26214, 26466, 26522, 26204, 25307, 23909, 23168, 22717, 22587, 
    22898, 23382, 24331, 25159, 26505, 26952, 27212, 26582, 26157, 25749, 
    24995, 24267,
  26171, 26163, 26473, 26513, 26247, 25271, 23991, 23171, 22651, 22642, 
    22963, 23439, 24236, 25323, 26531, 27019, 27334, 26724, 26168, 25685, 
    25078, 24360,
  26100, 26091, 26419, 26493, 26182, 25295, 23906, 23230, 22698, 22627, 
    22799, 23362, 24274, 25286, 26432, 26954, 27319, 26791, 26310, 25875, 
    25135, 24509,
  26057, 26055, 26357, 26390, 26150, 25229, 23955, 23194, 22730, 22626, 
    22860, 23418, 24070, 25275, 26414, 26868, 27288, 26687, 26301, 25840, 
    25295, 24589,
  26040, 26060, 26298, 26375, 26132, 25257, 23929, 23195, 22743, 22589, 
    22890, 23280, 24233, 25300, 26612, 26773, 27140, 26676, 26274, 25925, 
    25269, 24576,
  26008, 26057, 26338, 26382, 26145, 25240, 23971, 23233, 22751, 22617, 
    22879, 23409, 24290, 25518, 26434, 26754, 27079, 26655, 26224, 25820, 
    25231, 24709,
  25918, 26005, 26247, 26389, 26067, 25258, 23997, 23248, 22796, 22733, 
    22944, 23370, 24230, 25396, 26655, 26638, 27023, 26637, 26175, 25847, 
    25281, 24697,
  25775, 25894, 26182, 26319, 26074, 25257, 23967, 23254, 22771, 22630, 
    22834, 23288, 24147, 25422, 26593, 26517, 26932, 26491, 26182, 25710, 
    25293, 24683,
  25636, 25771, 26132, 26222, 26091, 25226, 23990, 23256, 22823, 22648, 
    22872, 23437, 24151, 25375, 26676, 26334, 26836, 26447, 26126, 25734, 
    25242, 24832,
  25556, 25677, 25915, 26117, 26000, 25223, 23969, 23254, 22796, 22722, 
    22900, 23391, 24002, 25452, 26457, 26170, 26866, 26453, 26147, 25809, 
    25357, 24852,
  25543, 25651, 26023, 26195, 26069, 25225, 24005, 23252, 22817, 22655, 
    22909, 23378, 24249, 25425, 26429, 26157, 26823, 26469, 26106, 25788, 
    25357, 24988,
  25570, 25677, 26101, 26217, 26082, 25233, 23983, 23285, 22826, 22694, 
    22949, 23398, 24215, 25199, 26554, 26156, 26729, 26386, 26016, 25707, 
    25313, 24916,
  25594, 25717, 26050, 26213, 26050, 25276, 24023, 23336, 22817, 22674, 
    22983, 23339, 24249, 25347, 26772, 26116, 26728, 26363, 26050, 25726, 
    25218, 24830,
  25618, 25755, 25997, 26220, 26056, 25290, 24025, 23319, 22842, 22674, 
    22953, 23339, 24221, 25455, 26288, 26005, 26875, 26463, 26001, 25658, 
    25245, 24831,
  25684, 25836, 25982, 26220, 26110, 25287, 24014, 23282, 22846, 22731, 
    22919, 23382, 24204, 25465, 26872, 25882, 26865, 26416, 25987, 25505, 
    25098, 24678,
  25819, 25978, 26136, 26337, 26178, 25292, 24006, 23300, 22840, 22613, 
    22873, 23401, 24308, 25395, 26668, 26006, 26829, 26356, 25872, 25505, 
    25042, 24531,
  25957, 26120, 26446, 26557, 26245, 25280, 24030, 23285, 22840, 22678, 
    22882, 23376, 24350, 25382, 26184, 26448, 26900, 26370, 25870, 25473, 
    24919, 24584,
  26007, 26170, 26563, 26632, 26264, 25354, 24034, 23284, 22880, 22721, 
    23015, 23411, 24212, 25172, 26401, 26678, 27104, 26382, 25847, 25369, 
    24856, 24424,
  25914, 26086, 26448, 26519, 26259, 25319, 24052, 23291, 22889, 22714, 
    22897, 23266, 24066, 25509, 26554, 26632, 27068, 26446, 25865, 25439, 
    24875, 24448,
  25741, 25929, 26200, 26325, 26154, 25287, 24015, 23329, 22893, 22718, 
    22854, 23388, 24375, 25248, 26413, 26315, 26896, 26441, 25832, 25334, 
    24816, 24446,
  25599, 25808, 26047, 26240, 26061, 25307, 23998, 23289, 22895, 22781, 
    22911, 23342, 24109, 25440, 26689, 26062, 26556, 26121, 25657, 25256, 
    24701, 24224,
  25582, 25792, 26162, 26291, 26125, 25281, 24040, 23323, 22880, 22685, 
    23019, 23370, 24066, 25438, 26524, 26203, 26479, 25988, 25531, 25204, 
    24721, 24277,
  25680, 25878, 26338, 26390, 26153, 25307, 24018, 23354, 22865, 22725, 
    22894, 23304, 24284, 25312, 26749, 26428, 26724, 26200, 25679, 25356, 
    24714, 24290,
  25824, 26015, 26469, 26447, 26187, 25318, 23986, 23307, 22897, 22720, 
    22930, 23343, 24374, 25244, 26751, 26626, 27090, 26491, 26015, 25483, 
    24834, 24311,
  25901, 26122, 26412, 26432, 26191, 25311, 24005, 23307, 22887, 22698, 
    22942, 23485, 24134, 25415, 26300, 26625, 27253, 26782, 26231, 25653, 
    24816, 24265,
  25829, 26094, 26325, 26333, 26112, 25301, 24028, 23338, 22907, 22749, 
    22938, 23375, 24242, 25454, 26866, 26511, 27224, 26819, 26269, 25656, 
    24847, 24298,
  25572, 25863, 26184, 26329, 26098, 25266, 24008, 23305, 22898, 22766, 
    22949, 23367, 24133, 25216, 26634, 26389, 27279, 26884, 26283, 25704, 
    24937, 24292,
  25101, 25388, 26075, 26263, 26107, 25246, 24014, 23309, 22860, 22778, 
    22939, 23352, 24426, 25331, 26841, 26278, 27187, 26875, 26313, 25729, 
    24962, 24339,
  24382, 24663, 25735, 26053, 26015, 25188, 23980, 23304, 22947, 22799, 
    23036, 23380, 24251, 25487, 26487, 25944, 27093, 26931, 26354, 25863, 
    25033, 24365,
  23413, 23713, 25245, 25737, 25891, 25170, 23978, 23260, 22901, 22765, 
    23000, 23358, 24152, 25457, 26495, 25310, 26846, 26950, 26492, 25869, 
    25185, 24534,
  22254, 22627, 24727, 25401, 25710, 25146, 23931, 23305, 22907, 22756, 
    22986, 23337, 24315, 25469, 26644, 24701, 26601, 26991, 26520, 25949, 
    25179, 24527,
  21057, 21522, 24143, 25047, 25537, 25087, 23949, 23317, 22905, 22824, 
    22945, 23412, 24104, 25358, 26333, 24206, 26501, 26866, 26415, 25864, 
    25150, 24481,
  20063, 20590, 23276, 24437, 25302, 24989, 23936, 23324, 22921, 22755, 
    23062, 23501, 24162, 25296, 26449, 23187, 25725, 26690, 26432, 25825, 
    25139, 24454,
  19493, 20035, 22657, 24068, 25115, 24942, 23957, 23271, 22929, 22814, 
    22992, 23408, 24325, 25365, 26469, 22376, 25249, 26716, 26434, 25964, 
    25191, 24503,
  19460, 19976, 22973, 24224, 25159, 24971, 23885, 23304, 22894, 22867, 
    23040, 23429, 24205, 25310, 26534, 22699, 25666, 26692, 26443, 25928, 
    25212, 24634,
  19895, 20343, 23534, 24544, 25256, 24937, 23906, 23307, 22970, 22817, 
    23004, 23494, 24281, 25383, 26555, 23295, 25860, 26734, 26477, 26003, 
    25270, 24650,
  20550, 20915, 23859, 24761, 25343, 24923, 23879, 23309, 22965, 22876, 
    22980, 23439, 24401, 25435, 26580, 23696, 25854, 26748, 26477, 25970, 
    25237, 24757,
  21150, 21450, 24024, 24951, 25411, 24962, 23879, 23325, 22939, 22855, 
    23029, 23417, 24344, 25563, 26787, 24006, 26040, 26784, 26411, 25996, 
    25315, 24690,
  21550, 21823, 24044, 24899, 25365, 24904, 23854, 23283, 23014, 22879, 
    23119, 23454, 24362, 25406, 26390, 24012, 25969, 26775, 26422, 25931, 
    25316, 24750,
  21750, 22028, 23994, 24868, 25378, 24959, 23854, 23272, 22966, 22909, 
    23048, 23501, 24207, 25337, 26769, 23930, 25907, 26699, 26338, 25941, 
    25233, 24652,
  21824, 22097, 23991, 24840, 25366, 24906, 23868, 23264, 22955, 22878, 
    23037, 23455, 24237, 25468, 26741, 23804, 25791, 26665, 26372, 25845, 
    25177, 24620,
  21827, 22055, 24079, 24864, 25358, 24857, 23821, 23289, 22949, 22929, 
    23111, 23571, 24404, 25470, 26601, 23898, 25767, 26575, 26238, 25805, 
    25159, 24641,
  21742, 21932, 24223, 24994, 25381, 24870, 23821, 23284, 22971, 22908, 
    23102, 23470, 24476, 25644, 27082, 24221, 26143, 26665, 26350, 25776, 
    25163, 24736,
  21572, 21774, 24248, 25013, 25385, 24867, 23768, 23263, 22942, 22893, 
    23141, 23495, 24358, 25437, 26778, 24443, 26266, 26641, 26337, 25723, 
    25239, 24694,
  21364, 21633, 23952, 24894, 25308, 24757, 23748, 23240, 22947, 22880, 
    23170, 23475, 24408, 25754, 26563, 24235, 26150, 26690, 26266, 25930, 
    25235, 24716,
  21203, 21533, 23711, 24762, 25289, 24772, 23731, 23248, 22974, 22861, 
    23109, 23608, 24450, 25484, 27038, 23952, 26062, 26571, 26245, 25884, 
    25262, 24703,
  21106, 21475, 23834, 24812, 25279, 24783, 23765, 23246, 22979, 22910, 
    23055, 23552, 24373, 25552, 26561, 23978, 26091, 26547, 26251, 25855, 
    25251, 24697,
  21015, 21398, 24065, 24956, 25326, 24708, 23731, 23235, 22942, 22904, 
    23167, 23518, 24430, 25668, 26693, 24253, 26184, 26524, 26100, 25744, 
    25187, 24572,
  20795, 21217, 24185, 25013, 25340, 24710, 23699, 23223, 22987, 22933, 
    23212, 23583, 24575, 25694, 26928, 24306, 26179, 26522, 26176, 25765, 
    25094, 24658,
  20395, 20854, 23857, 24848, 25324, 24729, 23694, 23210, 22987, 22928, 
    23091, 23551, 24439, 25704, 26736, 23960, 26124, 26563, 26167, 25754, 
    25178, 24693,
  19879, 20350, 23494, 24684, 25240, 24640, 23673, 23194, 23021, 22912, 
    23081, 23549, 24458, 25812, 26939, 23387, 26004, 26516, 26121, 25738, 
    25186, 24647,
  19479, 19869, 23304, 24585, 25167, 24621, 23639, 23186, 22992, 22993, 
    23176, 23643, 24432, 25462, 26582, 22979, 25797, 26482, 26095, 25640, 
    25124, 24521,
  19390, 19672, 23428, 24658, 25143, 24591, 23586, 23242, 22993, 22979, 
    23114, 23567, 24431, 25825, 26804, 22860, 25750, 26444, 26056, 25629, 
    25063, 24382,
  19731, 19895, 23449, 24668, 25220, 24592, 23599, 23204, 23047, 22947, 
    23209, 23604, 24664, 25980, 26925, 22826, 25640, 26368, 26051, 25670, 
    25076, 24410,
  20418, 20511, 23763, 24801, 25138, 24500, 23621, 23162, 23002, 22974, 
    23179, 23622, 24561, 25799, 26904, 23032, 25778, 26463, 26135, 25746, 
    25217, 24499,
  21249, 21318, 24273, 25048, 25243, 24523, 23556, 23149, 22949, 22955, 
    23219, 23643, 24692, 25822, 26941, 23732, 26031, 26520, 26205, 25875, 
    25243, 24687,
  21983, 22076, 24656, 25212, 25247, 24464, 23509, 23151, 23038, 22952, 
    23149, 23712, 24593, 25861, 26903, 24290, 26250, 26424, 26150, 25789, 
    25256, 24822,
  22498, 22612, 24759, 25330, 25293, 24458, 23462, 23175, 23020, 23055, 
    23159, 23682, 24523, 26113, 27104, 24453, 26132, 26373, 26079, 25776, 
    25140, 24669,
  22785, 22913, 24856, 25357, 25224, 24406, 23493, 23177, 23077, 23039, 
    23083, 23733, 24603, 25912, 26928, 24384, 26259, 26395, 26085, 25762, 
    25154, 24650,
  22941, 23079, 24964, 25402, 25229, 24388, 23441, 23167, 23040, 23029, 
    23240, 23737, 24595, 25845, 26884, 24369, 26236, 26396, 26007, 25848, 
    25118, 24570,
  23083, 23212, 25050, 25421, 25187, 24293, 23460, 23139, 23046, 23043, 
    23277, 23701, 24610, 25956, 27076, 24439, 26240, 26384, 26018, 25718, 
    25080, 24463,
  23278, 23366, 25155, 25458, 25199, 24290, 23438, 23132, 23076, 23089, 
    23290, 23801, 24729, 26184, 26889, 24549, 26241, 26274, 25950, 25651, 
    24992, 24463,
  23522, 23547, 25328, 25526, 25120, 24219, 23399, 23167, 23048, 23032, 
    23233, 23831, 24692, 25999, 27087, 24582, 26300, 26294, 25968, 25524, 
    24912, 24278,
  23762, 23754, 25408, 25572, 25112, 24162, 23398, 23177, 23059, 23005, 
    23268, 23811, 24868, 26103, 27229, 24687, 26246, 26275, 25890, 25490, 
    24965, 24287,
  23858, 23850, 25451, 25606, 25050, 24151, 23340, 23122, 23075, 23101, 
    23232, 23764, 24926, 26166, 27335, 24755, 26276, 26145, 25769, 25431, 
    24820, 24237,
  23710, 23681, 25545, 25590, 25001, 24012, 23333, 23121, 23112, 23082, 
    23340, 23898, 24793, 26137, 27028, 24926, 26271, 26078, 25639, 25217, 
    24658, 24165,
  23351, 23287, 25614, 25582, 24953, 23988, 23273, 23125, 23073, 23111, 
    23346, 23865, 24862, 26135, 27366, 24968, 26319, 26000, 25553, 25145, 
    24514, 24150,
  23171, 23068, 25635, 25536, 24865, 23920, 23244, 23129, 23082, 23084, 
    23259, 23879, 25011, 26355, 27087, 24905, 26309, 25904, 25540, 25110, 
    24489, 24031,
  27550, 27442, 27595, 27036, 25725, 24135, 22769, 22314, 22226, 22526, 
    22858, 23683, 24882, 25936, 26490, 28093, 27553, 26614, 26012, 25384, 
    24507, 23756,
  27524, 27416, 27493, 26982, 25796, 24222, 22807, 22370, 22214, 22484, 
    22925, 23522, 24655, 25654, 26596, 27826, 27126, 26358, 25847, 25278, 
    24462, 23816,
  27466, 27376, 27347, 26882, 25816, 24390, 22925, 22423, 22218, 22478, 
    22871, 23620, 24708, 25662, 26619, 27534, 26913, 26138, 25663, 25142, 
    24509, 23784,
  27371, 27329, 27210, 26810, 25888, 24467, 23015, 22415, 22269, 22519, 
    22976, 23576, 24598, 25597, 26871, 27391, 26969, 26092, 25569, 25079, 
    24477, 23770,
  27321, 27321, 27193, 26858, 25942, 24507, 23069, 22519, 22336, 22539, 
    22979, 23562, 24562, 25905, 26724, 27304, 26975, 26197, 25741, 25240, 
    24560, 23849,
  27267, 27281, 27063, 26786, 25953, 24579, 23130, 22545, 22294, 22525, 
    22961, 23562, 24632, 25750, 26806, 27108, 27073, 26301, 25812, 25253, 
    24585, 23915,
  27192, 27168, 26778, 26597, 25889, 24612, 23183, 22548, 22311, 22518, 
    22948, 23637, 24572, 25706, 26622, 26601, 26526, 26079, 25673, 25141, 
    24529, 23901,
  27510, 27366, 26700, 26375, 25713, 24549, 23237, 22498, 22266, 22479, 
    22882, 23364, 24463, 25631, 26557, 26198, 24984, 25175, 25093, 24844, 
    24340, 23848,
  27382, 27231, 26664, 26420, 25775, 24624, 23264, 22551, 22254, 22490, 
    22856, 23453, 24315, 25503, 26409, 26215, 24635, 24836, 24879, 24700, 
    24251, 23794,
  26830, 26810, 26653, 26527, 25959, 24728, 23353, 22672, 22406, 22508, 
    22896, 23388, 24410, 25567, 26823, 26488, 26226, 25747, 25471, 25004, 
    24433, 23915,
  26688, 26716, 26682, 26538, 25972, 24826, 23396, 22742, 22401, 22519, 
    22867, 23505, 24470, 25519, 26594, 26700, 26581, 25934, 25553, 25028, 
    24438, 23921,
  26602, 26654, 26689, 26556, 26040, 24804, 23482, 22757, 22445, 22567, 
    22834, 23443, 24371, 25676, 26579, 26732, 26379, 25945, 25537, 25013, 
    24493, 23893,
  26582, 26653, 26690, 26556, 26022, 24897, 23509, 22825, 22457, 22581, 
    22926, 23512, 24425, 25539, 26740, 26784, 26527, 26032, 25596, 25071, 
    24466, 23898,
  26639, 26714, 26718, 26597, 26113, 24978, 23523, 22842, 22412, 22571, 
    22895, 23477, 24389, 25834, 26596, 26965, 26941, 26280, 25737, 25100, 
    24477, 23843,
  26747, 26818, 26768, 26712, 26160, 24976, 23560, 22844, 22479, 22517, 
    22879, 23483, 24451, 25497, 26626, 27078, 26988, 26149, 25596, 25085, 
    24441, 23885,
  26866, 26912, 26860, 26737, 26191, 25085, 23610, 22908, 22493, 22636, 
    22867, 23445, 24256, 25647, 26951, 27096, 26676, 25916, 25525, 24989, 
    24415, 23849,
  26932, 26962, 26770, 26745, 26229, 25071, 23687, 22921, 22526, 22587, 
    22948, 23537, 24360, 25611, 26605, 27073, 26675, 26091, 25649, 25093, 
    24381, 23854,
  26913, 26950, 26763, 26679, 26204, 25040, 23660, 22959, 22537, 22522, 
    22811, 23381, 24267, 25429, 26666, 27048, 26955, 26391, 25862, 25317, 
    24576, 23919,
  26795, 26866, 26736, 26647, 26187, 25111, 23752, 22974, 22611, 22611, 
    22839, 23483, 24347, 25589, 26863, 26953, 26957, 26413, 25882, 25415, 
    24607, 23918,
  26603, 26685, 26614, 26590, 26134, 25068, 23735, 23029, 22575, 22578, 
    22850, 23449, 24303, 25529, 26474, 26831, 26644, 26284, 25910, 25438, 
    24646, 24126,
  26361, 26431, 26532, 26489, 26099, 25132, 23757, 23021, 22592, 22545, 
    22872, 23431, 24328, 25579, 26454, 26766, 26535, 26255, 25938, 25440, 
    24760, 24079,
  26115, 26169, 26444, 26457, 26132, 25112, 23736, 23024, 22585, 22576, 
    22932, 23437, 24367, 25375, 26744, 26768, 26543, 26282, 25903, 25453, 
    24854, 24139,
  25922, 25978, 26349, 26422, 26141, 25175, 23798, 23067, 22595, 22581, 
    22942, 23512, 24375, 25296, 26474, 26845, 26938, 26479, 26058, 25589, 
    24874, 24218,
  25820, 25903, 26438, 26465, 26166, 25196, 23807, 23086, 22618, 22531, 
    22870, 23383, 24246, 25540, 26766, 26899, 27057, 26633, 26150, 25737, 
    24994, 24317,
  25817, 25910, 26414, 26495, 26206, 25208, 23849, 23067, 22625, 22576, 
    22960, 23410, 24302, 25354, 26572, 26917, 27126, 26624, 26175, 25650, 
    24972, 24254,
  25874, 25945, 26325, 26474, 26179, 25207, 23830, 23145, 22653, 22590, 
    22884, 23332, 24216, 25421, 26678, 26922, 27141, 26650, 26209, 25716, 
    25053, 24406,
  25937, 25959, 26320, 26376, 26182, 25223, 23889, 23135, 22706, 22561, 
    22895, 23369, 24120, 25321, 26597, 26812, 27131, 26706, 26337, 25850, 
    25165, 24412,
  25968, 25950, 26222, 26396, 26195, 25198, 23916, 23143, 22717, 22626, 
    22923, 23393, 24229, 25231, 26818, 26710, 27075, 26663, 26266, 25741, 
    25095, 24437,
  25957, 25923, 26210, 26357, 26169, 25277, 23925, 23162, 22746, 22603, 
    22962, 23371, 24154, 25334, 26217, 26709, 27281, 26715, 26276, 25753, 
    25113, 24458,
  25925, 25898, 26207, 26418, 26213, 25244, 23941, 23147, 22769, 22655, 
    22876, 23436, 24273, 25289, 26699, 26716, 27322, 26682, 26322, 25889, 
    25310, 24619,
  25913, 25904, 26240, 26412, 26169, 25273, 23970, 23156, 22736, 22663, 
    22893, 23451, 24266, 25352, 26557, 26737, 27296, 26851, 26401, 25987, 
    25297, 24627,
  25967, 25985, 26210, 26360, 26128, 25242, 23953, 23190, 22771, 22672, 
    22881, 23403, 24215, 25190, 26673, 26706, 27201, 26741, 26400, 25963, 
    25317, 24815,
  26079, 26139, 26286, 26435, 26113, 25204, 23934, 23236, 22762, 22689, 
    22937, 23297, 24217, 25140, 26635, 26701, 26986, 26672, 26303, 25937, 
    25374, 24841,
  26200, 26304, 26467, 26439, 26116, 25246, 23954, 23221, 22712, 22670, 
    22900, 23339, 24284, 25336, 26506, 26759, 26893, 26592, 26266, 25901, 
    25406, 24808,
  26267, 26411, 26432, 26453, 26091, 25211, 23946, 23224, 22799, 22655, 
    22834, 23311, 24303, 25337, 26685, 26726, 26894, 26560, 26197, 25795, 
    25361, 24969,
  26255, 26425, 26545, 26464, 26154, 25240, 23969, 23203, 22792, 22673, 
    22898, 23353, 24082, 25334, 26259, 26692, 26878, 26508, 26066, 25803, 
    25360, 24827,
  26196, 26384, 26442, 26491, 26119, 25271, 23985, 23273, 22788, 22673, 
    22882, 23353, 24258, 25350, 26512, 26618, 26944, 26376, 26004, 25733, 
    25348, 24924,
  26148, 26334, 26422, 26459, 26126, 25257, 23995, 23271, 22855, 22656, 
    22921, 23411, 24185, 25339, 26548, 26535, 26904, 26456, 26038, 25801, 
    25379, 24957,
  26141, 26324, 26474, 26520, 26150, 25256, 23989, 23289, 22785, 22649, 
    22834, 23430, 24293, 25432, 26559, 26575, 26862, 26437, 26072, 25744, 
    25296, 24946,
  26171, 26350, 26540, 26459, 26157, 25222, 24019, 23293, 22820, 22642, 
    22876, 23420, 24212, 25346, 26594, 26597, 26781, 26316, 25956, 25626, 
    25170, 24840,
  26204, 26381, 26443, 26528, 26179, 25274, 23997, 23274, 22817, 22648, 
    23042, 23393, 24093, 25341, 26537, 26576, 26841, 26307, 25886, 25589, 
    25145, 24720,
  26226, 26396, 26454, 26554, 26157, 25257, 24000, 23269, 22839, 22665, 
    22906, 23447, 24225, 25484, 26494, 26459, 26876, 26213, 25795, 25408, 
    25000, 24554,
  26245, 26417, 26448, 26505, 26199, 25279, 24064, 23308, 22835, 22684, 
    22878, 23458, 24265, 25454, 26482, 26406, 26268, 25710, 25401, 25167, 
    24751, 24475,
  26262, 26438, 26636, 26607, 26208, 25318, 24018, 23309, 22885, 22713, 
    22891, 23386, 24340, 25517, 26861, 26496, 25716, 25203, 25059, 24850, 
    24548, 24300,
  26213, 26400, 26543, 26682, 26203, 25331, 24000, 23308, 22873, 22680, 
    22898, 23414, 24272, 25479, 26642, 26618, 26128, 25571, 25244, 24987, 
    24636, 24193,
  26051, 26245, 26482, 26507, 26220, 25296, 24035, 23331, 22860, 22720, 
    22916, 23326, 24142, 25548, 26619, 26578, 26290, 25735, 25399, 25050, 
    24598, 24233,
  25783, 25982, 26136, 26335, 26091, 25252, 24005, 23303, 22845, 22736, 
    22975, 23418, 24302, 25461, 26437, 26299, 26515, 26073, 25610, 25158, 
    24681, 24385,
  25523, 25716, 26031, 26206, 26106, 25279, 23986, 23290, 22858, 22762, 
    23057, 23415, 24214, 25550, 26704, 26062, 26455, 26060, 25571, 25221, 
    24673, 24215,
  25382, 25572, 25910, 26150, 26056, 25254, 24024, 23325, 22863, 22746, 
    23009, 23420, 24202, 25381, 26649, 25837, 26371, 26109, 25576, 25168, 
    24692, 24221,
  25424, 25609, 25921, 26179, 26057, 25279, 24003, 23323, 22910, 22773, 
    23051, 23423, 24272, 25117, 26886, 25987, 26612, 26294, 25816, 25259, 
    24788, 24240,
  25600, 25786, 26190, 26397, 26182, 25290, 24030, 23337, 22874, 22739, 
    22946, 23390, 24347, 25604, 27121, 26353, 26987, 26520, 26067, 25479, 
    24870, 24287,
  25814, 26004, 26451, 26535, 26214, 25279, 24008, 23298, 22903, 22765, 
    22946, 23385, 24269, 25583, 26491, 26670, 27328, 26768, 26216, 25662, 
    24958, 24476,
  25943, 26152, 26500, 26547, 26216, 25314, 24045, 23322, 22909, 22772, 
    22940, 23392, 24256, 25549, 26632, 26729, 27454, 26871, 26316, 25708, 
    25042, 24523,
  25898, 26125, 26329, 26500, 26196, 25316, 24019, 23296, 22892, 22798, 
    23033, 23494, 24379, 25498, 26846, 26601, 27419, 26924, 26340, 25834, 
    25036, 24476,
  25635, 25878, 26200, 26375, 26101, 25308, 23999, 23329, 22913, 22773, 
    22990, 23460, 24284, 25454, 26638, 26400, 27194, 26894, 26347, 25903, 
    25125, 24658,
  25115, 25378, 26070, 26265, 26101, 25246, 23984, 23326, 22904, 22774, 
    23097, 23481, 24302, 25441, 26550, 26287, 27238, 26963, 26468, 25854, 
    25189, 24570,
  24312, 24614, 25940, 26182, 26041, 25273, 24017, 23312, 22974, 22802, 
    23006, 23374, 24319, 25527, 26425, 26090, 27250, 27012, 26521, 25862, 
    25201, 24705,
  23262, 23618, 25448, 25845, 25926, 25195, 23962, 23265, 22889, 22819, 
    22950, 23440, 24415, 25387, 26972, 25575, 27072, 27010, 26479, 25999, 
    25271, 24625,
  22082, 22519, 24623, 25337, 25642, 25127, 23985, 23301, 22925, 22819, 
    23064, 23445, 24097, 25413, 26565, 24782, 26572, 26842, 26432, 25892, 
    25228, 24592,
  20967, 21474, 23853, 24795, 25444, 25051, 23937, 23263, 22952, 22806, 
    23046, 23496, 24406, 25438, 26477, 23820, 26104, 26731, 26403, 25962, 
    25281, 24592,
  20153, 20681, 23045, 24358, 25178, 24995, 23928, 23332, 22921, 22866, 
    23021, 23390, 24285, 25402, 26794, 22879, 25459, 26743, 26482, 25924, 
    25168, 24532,
  19793, 20301, 22847, 24169, 25156, 24985, 23921, 23330, 22926, 22905, 
    23053, 23462, 24408, 25441, 26272, 22486, 25312, 26638, 26449, 25938, 
    25341, 24654,
  19921, 20386, 23168, 24363, 25241, 24979, 23898, 23315, 22952, 22884, 
    23039, 23509, 24251, 25334, 27082, 22950, 25594, 26738, 26500, 26082, 
    25310, 24699,
  20417, 20812, 23683, 24622, 25335, 24932, 23879, 23265, 22988, 22842, 
    23036, 23592, 24318, 25265, 26588, 23544, 25849, 26743, 26471, 26014, 
    25387, 24681,
  21032, 21351, 24047, 24878, 25362, 24983, 23954, 23296, 22921, 22915, 
    23087, 23557, 24318, 25529, 26931, 24017, 26073, 26772, 26486, 26013, 
    25393, 24768,
  21530, 21793, 24082, 24899, 25386, 24929, 23867, 23321, 22921, 22886, 
    23158, 23513, 24409, 25766, 26912, 24054, 25997, 26721, 26496, 26057, 
    25439, 24915,
  21816, 22059, 24010, 24857, 25360, 24943, 23897, 23297, 22956, 22926, 
    23066, 23536, 24430, 25734, 26678, 23851, 25722, 26727, 26450, 25994, 
    25300, 24754,
  21920, 22165, 24052, 24840, 25374, 24906, 23835, 23269, 22928, 22968, 
    23106, 23584, 24261, 25373, 26568, 23875, 25803, 26651, 26306, 25847, 
    25275, 24784,
  21916, 22147, 24033, 24868, 25356, 24929, 23824, 23288, 23005, 22917, 
    23135, 23594, 24381, 25641, 26759, 23839, 25806, 26646, 26325, 25844, 
    25225, 24718,
  21834, 22023, 24121, 24915, 25353, 24830, 23816, 23250, 22961, 22937, 
    23067, 23487, 24369, 25530, 26826, 24010, 25986, 26606, 26281, 25847, 
    25188, 24693,
  21643, 21816, 24200, 24982, 25379, 24818, 23828, 23264, 22994, 22933, 
    23186, 23470, 24369, 25563, 26688, 24336, 26213, 26638, 26303, 25818, 
    25223, 24707,
  21363, 21570, 23903, 24812, 25275, 24778, 23742, 23239, 22957, 22950, 
    23136, 23458, 24450, 25538, 26999, 24227, 26136, 26630, 26256, 25778, 
    25268, 24791,
  21081, 21358, 23589, 24640, 25248, 24751, 23723, 23243, 22932, 22937, 
    23149, 23581, 24436, 25635, 26754, 23812, 25928, 26635, 26254, 25823, 
    25237, 24861,
  20927, 21247, 23442, 24570, 25221, 24756, 23730, 23227, 22957, 22920, 
    23150, 23564, 24435, 25734, 26799, 23682, 25839, 26560, 26260, 25838, 
    25316, 24781,
  20941, 21277, 23654, 24653, 25237, 24730, 23733, 23232, 22985, 22962, 
    23153, 23658, 24404, 25596, 26676, 23834, 25912, 26550, 26198, 25829, 
    25325, 24801,
  21052, 21392, 24025, 24909, 25332, 24698, 23750, 23203, 22980, 22982, 
    23131, 23553, 24522, 25567, 26706, 24240, 26167, 26512, 26213, 25743, 
    25274, 24844,
  21084, 21477, 24190, 24988, 25342, 24663, 23701, 23202, 22966, 22960, 
    23142, 23696, 24500, 25783, 26828, 24469, 26355, 26568, 26178, 25858, 
    25326, 24696,
  20946, 21400, 24184, 24962, 25283, 24712, 23678, 23244, 23015, 23031, 
    23197, 23706, 24297, 25763, 26875, 24337, 26294, 26565, 26162, 25754, 
    25257, 24737,
  20661, 21145, 23887, 24883, 25281, 24669, 23661, 23235, 22990, 22994, 
    23236, 23650, 24548, 25636, 26952, 23893, 26100, 26526, 26178, 25750, 
    25260, 24658,
  20411, 20822, 23843, 24848, 25237, 24613, 23673, 23207, 22983, 23061, 
    23117, 23741, 24462, 25847, 27023, 23643, 25824, 26463, 26075, 25744, 
    25134, 24472,
  20346, 20651, 23942, 24899, 25215, 24597, 23632, 23215, 23008, 23053, 
    23173, 23696, 24595, 25716, 26662, 23621, 25994, 26484, 26092, 25765, 
    25098, 24520,
  20564, 20756, 24055, 24928, 25237, 24531, 23604, 23192, 23033, 23040, 
    23268, 23705, 24575, 25769, 27006, 23558, 25934, 26501, 26184, 25806, 
    25194, 24622,
  21016, 21142, 24146, 25034, 25276, 24557, 23582, 23182, 22997, 23062, 
    23171, 23802, 24641, 25963, 27129, 23624, 25966, 26496, 26172, 25801, 
    25290, 24670,
  21578, 21681, 24430, 25141, 25253, 24549, 23548, 23231, 23057, 23075, 
    23331, 23582, 24679, 26100, 26759, 23978, 26144, 26458, 26220, 25918, 
    25284, 24751,
  22091, 22219, 24676, 25266, 25268, 24509, 23542, 23200, 23012, 23049, 
    23213, 23660, 24668, 25951, 27038, 24278, 26194, 26470, 26187, 25831, 
    25348, 24753,
  22482, 22635, 24744, 25321, 25295, 24430, 23507, 23198, 23061, 23037, 
    23279, 23717, 24621, 25835, 27201, 24325, 26022, 26491, 26199, 25831, 
    25240, 24734,
  22738, 22911, 24848, 25321, 25202, 24404, 23501, 23182, 23053, 23115, 
    23178, 23717, 24850, 26190, 26744, 24337, 26131, 26448, 26135, 25811, 
    25201, 24694,
  22921, 23102, 24898, 25423, 25181, 24369, 23468, 23193, 23075, 23037, 
    23236, 23661, 24547, 25925, 27199, 24384, 26187, 26391, 26038, 25679, 
    25185, 24641,
  23106, 23267, 25050, 25479, 25206, 24308, 23451, 23203, 23070, 23096, 
    23224, 23756, 24769, 26091, 27288, 24453, 26211, 26481, 26094, 25641, 
    25115, 24474,
  23337, 23446, 25160, 25462, 25131, 24326, 23436, 23191, 23057, 23085, 
    23252, 23743, 24849, 26046, 27084, 24533, 26250, 26319, 25979, 25662, 
    25116, 24555,
  23608, 23644, 25289, 25525, 25106, 24206, 23390, 23143, 23098, 23100, 
    23291, 23841, 24759, 26044, 27179, 24605, 26340, 26325, 26018, 25566, 
    25042, 24515,
  23872, 23862, 25416, 25585, 25069, 24171, 23351, 23165, 23059, 23162, 
    23283, 23859, 24830, 26181, 27401, 24671, 26222, 26241, 25946, 25421, 
    24956, 24404,
  23985, 23970, 25451, 25565, 25074, 24115, 23372, 23175, 23128, 23068, 
    23265, 23801, 24937, 26097, 27242, 24795, 26228, 26262, 25888, 25405, 
    24906, 24374,
  23847, 23824, 25565, 25584, 25048, 24040, 23341, 23137, 23090, 23058, 
    23332, 23857, 24910, 26169, 27383, 24965, 26186, 26051, 25717, 25310, 
    24737, 24210,
  23492, 23457, 25571, 25573, 24985, 24005, 23296, 23186, 23137, 23087, 
    23333, 23897, 24816, 26163, 26848, 25055, 26333, 26053, 25629, 25132, 
    24619, 24133,
  23312, 23252, 25580, 25500, 24884, 23954, 23270, 23129, 23064, 23080, 
    23257, 24033, 24923, 26328, 27371, 24970, 26329, 25957, 25520, 25034, 
    24581, 24048,
  27461, 27384, 27500, 26932, 25723, 24157, 22789, 22346, 22207, 22531, 
    22931, 23682, 24576, 25844, 26532, 27943, 27466, 26429, 25844, 25240, 
    24359, 23607,
  27434, 27354, 27363, 26853, 25822, 24225, 22858, 22349, 22224, 22593, 
    22956, 23652, 24815, 25928, 27119, 27607, 27102, 26210, 25701, 25115, 
    24448, 23787,
  27375, 27305, 27257, 26728, 25759, 24305, 22945, 22437, 22211, 22627, 
    22992, 23696, 24713, 25734, 26853, 27313, 26832, 26134, 25647, 25135, 
    24513, 23935,
  27285, 27255, 27072, 26709, 25800, 24432, 23003, 22449, 22273, 22596, 
    22940, 23634, 24393, 26022, 26738, 27167, 26877, 26189, 25733, 25189, 
    24539, 24054,
  27245, 27256, 27000, 26683, 25826, 24470, 23057, 22515, 22284, 22550, 
    22985, 23593, 24722, 25632, 27149, 26929, 26907, 26259, 25781, 25337, 
    24582, 23980,
  27206, 27237, 26850, 26622, 25843, 24548, 23136, 22538, 22307, 22573, 
    22935, 23614, 24563, 25623, 26822, 26629, 26370, 25908, 25596, 25184, 
    24539, 23920,
  27572, 27497, 26751, 26428, 25728, 24526, 23138, 22497, 22241, 22496, 
    22905, 23543, 24611, 25765, 27116, 26418, 25575, 25539, 25277, 24992, 
    24390, 23900,
  27520, 27388, 26789, 26445, 25782, 24613, 23187, 22517, 22297, 22501, 
    22842, 23507, 24473, 25523, 26847, 26356, 24803, 25041, 25070, 24799, 
    24326, 23866,
  27439, 27290, 26840, 26544, 25799, 24658, 23273, 22538, 22270, 22495, 
    22862, 23550, 24487, 25657, 26560, 26635, 25649, 25423, 25180, 24823, 
    24364, 23866,
  26918, 26896, 26804, 26657, 25985, 24714, 23345, 22698, 22343, 22533, 
    22929, 23581, 24573, 25561, 26938, 26844, 26631, 25994, 25498, 25053, 
    24367, 23900,
  26778, 26812, 26779, 26649, 26035, 24739, 23419, 22715, 22426, 22639, 
    22935, 23467, 24439, 25701, 26312, 26965, 26669, 25901, 25440, 24959, 
    24335, 23926,
  26662, 26736, 26772, 26639, 26034, 24856, 23465, 22760, 22432, 22610, 
    22948, 23559, 24533, 25642, 26803, 26960, 26641, 25955, 25528, 25024, 
    24498, 23931,
  26597, 26698, 26703, 26634, 26049, 24891, 23476, 22839, 22482, 22624, 
    22837, 23532, 24447, 25607, 26732, 26970, 26826, 26085, 25613, 25070, 
    24426, 23923,
  26612, 26713, 26696, 26640, 26109, 24978, 23556, 22841, 22474, 22542, 
    22962, 23434, 24320, 25676, 26575, 27032, 27165, 26341, 25790, 25242, 
    24557, 24068,
  26693, 26780, 26713, 26688, 26115, 25001, 23562, 22855, 22489, 22573, 
    22859, 23401, 24465, 25722, 26887, 27106, 27200, 26490, 25869, 25308, 
    24573, 23943,
  26802, 26859, 26741, 26675, 26101, 25000, 23602, 22898, 22529, 22632, 
    22895, 23453, 24303, 25687, 26711, 27109, 27200, 26532, 25992, 25323, 
    24559, 23854,
  26866, 26917, 26821, 26699, 26199, 25023, 23665, 22950, 22587, 22612, 
    23002, 23531, 24444, 25521, 26531, 27044, 27211, 26506, 26004, 25365, 
    24595, 24000,
  26851, 26920, 26740, 26666, 26115, 25029, 23662, 22958, 22551, 22614, 
    22833, 23418, 24423, 25572, 26491, 27005, 27093, 26546, 26122, 25464, 
    24587, 24017,
  26737, 26840, 26580, 26601, 26132, 25068, 23720, 22970, 22562, 22597, 
    22936, 23448, 24282, 25592, 26500, 26852, 26938, 26525, 26053, 25537, 
    24701, 23915,
  26547, 26648, 26587, 26590, 26118, 25092, 23717, 23001, 22591, 22592, 
    22890, 23531, 24409, 25425, 26788, 26721, 26626, 26316, 25970, 25530, 
    24759, 24144,
  26302, 26378, 26500, 26492, 26115, 25118, 23776, 23047, 22623, 22603, 
    22911, 23479, 24321, 25343, 26499, 26691, 26604, 26266, 25881, 25495, 
    24840, 24144,
  26062, 26109, 26413, 26449, 26128, 25128, 23737, 23035, 22619, 22590, 
    22855, 23453, 24258, 25421, 26893, 26737, 26724, 26351, 26019, 25577, 
    24803, 24224,
  25885, 25929, 26411, 26451, 26148, 25187, 23853, 23099, 22693, 22664, 
    22932, 23446, 24404, 25490, 26584, 26825, 26938, 26525, 26091, 25625, 
    24917, 24256,
  25799, 25877, 26393, 26467, 26170, 25167, 23844, 23083, 22704, 22597, 
    22873, 23480, 24299, 25331, 26297, 26854, 26997, 26614, 26210, 25722, 
    24973, 24435,
  25795, 25901, 26309, 26482, 26181, 25145, 23831, 23112, 22637, 22660, 
    22843, 23514, 24290, 25418, 26791, 26894, 27127, 26684, 26222, 25760, 
    25065, 24320,
  25828, 25927, 26316, 26444, 26140, 25199, 23874, 23153, 22661, 22693, 
    22979, 23457, 24426, 25373, 26734, 26865, 27286, 26725, 26284, 25864, 
    25166, 24424,
  25851, 25897, 26260, 26412, 26154, 25222, 23906, 23164, 22696, 22621, 
    22840, 23514, 24200, 25546, 26445, 26678, 26895, 26572, 26266, 25743, 
    25037, 24497,
  25840, 25827, 26204, 26380, 26165, 25226, 23912, 23171, 22748, 22635, 
    22985, 23393, 24251, 25441, 26824, 26610, 26814, 26449, 26097, 25654, 
    25011, 24410,
  25800, 25752, 26131, 26415, 26154, 25271, 23920, 23167, 22748, 22649, 
    22950, 23466, 24292, 25210, 26764, 26622, 27271, 26740, 26357, 25901, 
    25226, 24583,
  25759, 25715, 26190, 26369, 26207, 25280, 23922, 23226, 22779, 22644, 
    22933, 23439, 24381, 25436, 26684, 26690, 27287, 26816, 26429, 25982, 
    25360, 24811,
  25765, 25748, 26194, 26361, 26141, 25311, 23958, 23241, 22790, 22678, 
    22842, 23528, 24335, 25271, 26168, 26643, 27179, 26775, 26391, 25953, 
    25385, 24927,
  25866, 25893, 26193, 26304, 26124, 25254, 23994, 23234, 22808, 22663, 
    22876, 23421, 24234, 25433, 26322, 26603, 27148, 26693, 26383, 25987, 
    25462, 24907,
  26062, 26148, 26363, 26363, 26091, 25215, 23964, 23253, 22795, 22617, 
    22903, 23430, 24330, 25332, 26565, 26664, 26943, 26488, 26266, 25922, 
    25507, 24987,
  26305, 26445, 26501, 26424, 26115, 25197, 23992, 23221, 22844, 22682, 
    22954, 23436, 24129, 25429, 26663, 26740, 26838, 26516, 26237, 25862, 
    25500, 25040,
  26514, 26693, 26540, 26472, 26150, 25199, 23963, 23250, 22815, 22681, 
    22826, 23446, 24322, 25562, 26627, 26744, 26776, 26447, 26147, 25695, 
    25423, 25048,
  26628, 26831, 26597, 26502, 26153, 25240, 23946, 23244, 22870, 22698, 
    22878, 23381, 24254, 25453, 26403, 26756, 26810, 26367, 26079, 25682, 
    25359, 25027,
  26651, 26879, 26648, 26556, 26149, 25248, 23973, 23269, 22789, 22724, 
    22978, 23391, 24219, 25167, 26498, 26801, 26814, 26344, 26003, 25639, 
    25186, 24935,
  26638, 26877, 26703, 26616, 26159, 25285, 23987, 23306, 22863, 22678, 
    22870, 23475, 24146, 25493, 26734, 26801, 26900, 26357, 25932, 25433, 
    25123, 24774,
  26636, 26876, 26704, 26635, 26182, 25272, 24019, 23289, 22833, 22720, 
    22962, 23461, 24150, 25438, 26431, 26784, 26938, 26375, 25932, 25507, 
    25110, 24722,
  26661, 26882, 26699, 26591, 26209, 25306, 24039, 23328, 22901, 22673, 
    22890, 23421, 24086, 25508, 26404, 26783, 26826, 26218, 25844, 25401, 
    24989, 24597,
  26678, 26873, 26604, 26653, 26251, 25287, 24020, 23279, 22895, 22728, 
    22936, 23468, 24226, 25451, 26822, 26731, 26794, 26138, 25698, 25363, 
    24946, 24517,
  26654, 26825, 26660, 26648, 26261, 25290, 24037, 23306, 22873, 22745, 
    22872, 23374, 24228, 25234, 26596, 26695, 25979, 25539, 25386, 25083, 
    24698, 24338,
  26570, 26739, 26629, 26624, 26269, 25309, 24053, 23319, 22882, 22687, 
    22869, 23395, 24206, 25448, 26360, 26571, 25434, 25071, 24992, 24911, 
    24558, 24218,
  26413, 26596, 26657, 26656, 26251, 25354, 24010, 23340, 22834, 22739, 
    22883, 23399, 24278, 25395, 26519, 26606, 25654, 25271, 25085, 24849, 
    24565, 24151,
  26146, 26354, 26603, 26610, 26236, 25294, 24017, 23337, 22898, 22746, 
    22951, 23356, 24210, 25415, 26356, 26628, 26384, 25863, 25573, 25079, 
    24660, 24224,
  25779, 26004, 26324, 26402, 26179, 25334, 24034, 23336, 22908, 22731, 
    22918, 23370, 24282, 25381, 26673, 26379, 26041, 25551, 25232, 24955, 
    24616, 24237,
  25377, 25604, 26018, 26231, 26037, 25289, 24001, 23341, 22847, 22793, 
    22924, 23451, 24327, 25332, 26411, 26033, 25887, 25535, 25271, 24858, 
    24597, 24148,
  25070, 25277, 25853, 26143, 26018, 25273, 24015, 23337, 22927, 22826, 
    23029, 23436, 24235, 25404, 26741, 25878, 26431, 25956, 25584, 25145, 
    24665, 24160,
  24953, 25141, 25825, 26128, 26000, 25240, 24012, 23309, 22914, 22768, 
    22958, 23367, 24177, 25565, 26635, 25806, 26809, 26459, 25953, 25490, 
    24856, 24300,
  25045, 25228, 25815, 26104, 26052, 25295, 24001, 23351, 22878, 22831, 
    22935, 23411, 24174, 25321, 26868, 25816, 26825, 26659, 26145, 25569, 
    24900, 24426,
  25262, 25463, 26049, 26236, 26114, 25293, 24025, 23339, 22905, 22782, 
    22917, 23426, 24137, 25445, 26624, 26194, 27044, 26760, 26196, 25671, 
    25002, 24386,
  25493, 25710, 26372, 26481, 26232, 25315, 24010, 23327, 22872, 22822, 
    22965, 23456, 24111, 25291, 26363, 26625, 27435, 26938, 26304, 25729, 
    24950, 24426,
  25616, 25837, 26554, 26547, 26268, 25330, 24023, 23324, 22910, 22769, 
    23020, 23461, 24294, 25390, 26375, 26786, 27554, 26896, 26307, 25756, 
    25015, 24487,
  25543, 25753, 26418, 26476, 26168, 25315, 24018, 23337, 22949, 22760, 
    22936, 23411, 24404, 25354, 26784, 26678, 27438, 26954, 26379, 25851, 
    25002, 24481,
  25235, 25451, 26213, 26326, 26109, 25313, 24015, 23363, 22929, 22739, 
    23058, 23400, 24237, 25317, 26563, 26436, 27275, 26984, 26421, 25871, 
    25187, 24623,
  24669, 24926, 26042, 26265, 26086, 25251, 23994, 23326, 22940, 22832, 
    22963, 23426, 24336, 25396, 26428, 26281, 27294, 26996, 26500, 25921, 
    25181, 24515,
  23851, 24179, 25777, 26034, 25978, 25242, 23977, 23314, 22934, 22761, 
    22908, 23329, 24334, 25442, 26613, 26119, 27251, 26979, 26457, 25922, 
    25193, 24595,
  22849, 23244, 25319, 25775, 25804, 25124, 23957, 23285, 22944, 22824, 
    22950, 23390, 24142, 25420, 25987, 25647, 27117, 26882, 26463, 25849, 
    25168, 24489,
  21799, 22260, 24406, 25142, 25565, 25062, 23931, 23322, 22935, 22810, 
    22954, 23448, 24265, 25398, 26683, 24599, 26659, 26809, 26429, 25916, 
    25187, 24429,
  20891, 21387, 23590, 24615, 25361, 25031, 23939, 23307, 22898, 22855, 
    22909, 23499, 24211, 25278, 26277, 23518, 25856, 26690, 26387, 25879, 
    25145, 24610,
  20316, 20799, 23301, 24425, 25247, 24994, 23930, 23338, 22928, 22883, 
    23049, 23362, 24339, 25342, 26404, 23094, 25790, 26653, 26419, 25966, 
    25307, 24651,
  20161, 20606, 23497, 24474, 25262, 24936, 23927, 23326, 22975, 22833, 
    23037, 23481, 24272, 25314, 26510, 23095, 25718, 26722, 26460, 26018, 
    25352, 24666,
  20398, 20805, 23607, 24609, 25304, 24993, 23904, 23292, 22928, 22818, 
    22984, 23500, 24293, 25570, 26597, 23485, 25906, 26741, 26512, 25981, 
    25334, 24764,
  20895, 21246, 23872, 24772, 25355, 24914, 23907, 23271, 22910, 22860, 
    23056, 23402, 24058, 25393, 26538, 23803, 25993, 26703, 26442, 26019, 
    25412, 24865,
  21435, 21721, 24139, 24917, 25389, 24960, 23890, 23281, 22931, 22846, 
    23067, 23443, 24343, 25506, 26640, 24059, 26061, 26725, 26415, 26029, 
    25418, 24785,
  21834, 22069, 24149, 24959, 25336, 24906, 23849, 23248, 22929, 22915, 
    23044, 23483, 24360, 25625, 26191, 24023, 25923, 26644, 26431, 25943, 
    25310, 24726,
  22033, 22249, 24062, 24930, 25330, 24904, 23865, 23276, 22946, 22893, 
    23097, 23499, 24299, 25679, 26660, 23890, 25809, 26572, 26346, 25910, 
    25330, 24752,
  22071, 22290, 24068, 24875, 25300, 24857, 23843, 23237, 22921, 22854, 
    23024, 23476, 24404, 25451, 26414, 23872, 25928, 26553, 26290, 25814, 
    25223, 24742,
  22007, 22215, 24032, 24912, 25337, 24813, 23778, 23219, 22910, 22917, 
    23126, 23534, 24386, 25501, 26451, 23876, 25843, 26626, 26330, 25886, 
    25204, 24676,
  21850, 22029, 24160, 24944, 25328, 24863, 23752, 23226, 22971, 22876, 
    23200, 23441, 24485, 25346, 26985, 24130, 26098, 26572, 26334, 25784, 
    25327, 24878,
  21566, 21744, 24041, 24907, 25308, 24842, 23764, 23269, 22984, 22850, 
    23126, 23493, 24436, 25648, 26809, 24235, 26238, 26671, 26349, 25829, 
    25298, 24853,
  21192, 21409, 23694, 24662, 25236, 24769, 23748, 23280, 22985, 22898, 
    23142, 23583, 24374, 25483, 26367, 23836, 26056, 26633, 26296, 25864, 
    25343, 24817,
  20849, 21122, 23349, 24476, 25206, 24807, 23777, 23290, 22989, 22893, 
    23057, 23635, 24295, 25597, 26570, 23478, 25766, 26616, 26328, 25797, 
    25415, 24879,
  20697, 20990, 23346, 24530, 25204, 24769, 23749, 23264, 22976, 22961, 
    23044, 23628, 24451, 25448, 26873, 23490, 25896, 26476, 26224, 25850, 
    25308, 24792,
  20791, 21079, 23675, 24665, 25252, 24730, 23735, 23299, 22995, 22979, 
    23173, 23636, 24422, 25664, 26609, 23756, 26031, 26453, 26217, 25809, 
    25323, 24753,
  21051, 21333, 23982, 24864, 25287, 24741, 23714, 23257, 23002, 22993, 
    23117, 23614, 24483, 25584, 27001, 24178, 26149, 26530, 26245, 25741, 
    25182, 24682,
  21279, 21614, 24280, 24994, 25282, 24690, 23689, 23242, 23003, 23009, 
    23130, 23585, 24453, 25730, 26650, 24468, 26349, 26484, 26162, 25676, 
    25223, 24754,
  21356, 21763, 24294, 25054, 25315, 24670, 23705, 23223, 23042, 23012, 
    23149, 23671, 24497, 25847, 26854, 24463, 26294, 26482, 26139, 25728, 
    25097, 24668,
  21271, 21728, 24240, 25061, 25331, 24668, 23679, 23222, 23035, 23026, 
    23137, 23536, 24573, 25757, 27482, 24295, 26218, 26486, 26126, 25668, 
    25131, 24522,
  21161, 21570, 24235, 25031, 25292, 24668, 23651, 23247, 23043, 22993, 
    23103, 23635, 24509, 25812, 26982, 24158, 26154, 26494, 26101, 25626, 
    25030, 24570,
  21133, 21464, 24285, 25042, 25264, 24597, 23611, 23206, 23012, 22973, 
    23067, 23683, 24607, 25819, 27097, 24107, 26081, 26479, 26125, 25728, 
    25058, 24565,
  21263, 21506, 24299, 25068, 25285, 24578, 23593, 23192, 23046, 23023, 
    23276, 23680, 24762, 25937, 26884, 24045, 26015, 26475, 26203, 25685, 
    25237, 24753,
  21526, 21714, 24360, 25139, 25248, 24540, 23570, 23252, 23042, 23048, 
    23197, 23665, 24530, 25982, 26776, 23992, 26066, 26499, 26183, 25812, 
    25232, 24722,
  21861, 22017, 24442, 25190, 25239, 24503, 23533, 23201, 23041, 23097, 
    23183, 23699, 24583, 25882, 26881, 24081, 26046, 26396, 26163, 25724, 
    25232, 24756,
  22179, 22342, 24601, 25218, 25257, 24483, 23527, 23185, 23036, 23057, 
    23252, 23724, 24559, 25762, 27104, 24190, 26071, 26473, 26143, 25805, 
    25251, 24791,
  22458, 22630, 24674, 25275, 25273, 24441, 23542, 23215, 23039, 23074, 
    23342, 23694, 24594, 25944, 26788, 24236, 26109, 26437, 26121, 25774, 
    25194, 24605,
  22691, 22869, 24796, 25340, 25240, 24398, 23500, 23176, 23101, 23078, 
    23158, 23842, 24623, 25941, 27191, 24309, 26150, 26386, 26043, 25697, 
    25245, 24645,
  22909, 23082, 24955, 25401, 25242, 24357, 23498, 23201, 23085, 23079, 
    23269, 23762, 24542, 25812, 27109, 24400, 26226, 26336, 26049, 25678, 
    25119, 24585,
  23145, 23292, 25106, 25498, 25198, 24335, 23482, 23226, 23056, 23043, 
    23244, 23709, 24688, 25934, 27109, 24451, 26248, 26368, 25996, 25566, 
    25043, 24566,
  23412, 23514, 25255, 25503, 25194, 24229, 23445, 23178, 23085, 23091, 
    23248, 23749, 24701, 25924, 26950, 24550, 26200, 26338, 25976, 25568, 
    25102, 24512,
  23699, 23739, 25354, 25490, 25142, 24214, 23399, 23222, 23120, 23071, 
    23290, 23844, 24789, 25938, 26644, 24535, 26147, 26292, 25906, 25503, 
    24983, 24440,
  23966, 23961, 25361, 25566, 25104, 24159, 23349, 23188, 23108, 23116, 
    23255, 23852, 24775, 26084, 27032, 24601, 26167, 26229, 25819, 25482, 
    24954, 24349,
  24080, 24060, 25434, 25530, 25012, 24117, 23351, 23210, 23079, 23063, 
    23276, 23883, 24725, 25937, 27007, 24731, 26185, 26107, 25755, 25423, 
    24828, 24292,
  23944, 23915, 25536, 25584, 24943, 24014, 23326, 23131, 23106, 23075, 
    23244, 23941, 24792, 26153, 27314, 24893, 26187, 25997, 25679, 25295, 
    24723, 24128,
  23592, 23565, 25572, 25530, 24914, 24021, 23295, 23171, 23101, 23070, 
    23301, 23926, 24976, 26226, 27186, 25033, 26302, 25956, 25573, 25149, 
    24618, 24037,
  23414, 23371, 25606, 25506, 24887, 23945, 23256, 23175, 23084, 23197, 
    23307, 23945, 24970, 26251, 27428, 24998, 26304, 25924, 25456, 25007, 
    24446, 23892,
  27387, 27344, 27403, 26891, 25712, 24120, 22754, 22345, 22268, 22555, 
    22917, 23717, 24750, 25977, 26553, 27796, 27338, 26395, 25797, 25135, 
    24287, 23645,
  27362, 27314, 27263, 26872, 25751, 24227, 22854, 22339, 22241, 22594, 
    22905, 23637, 24653, 25635, 26894, 27606, 27173, 26190, 25653, 25146, 
    24479, 23858,
  27311, 27266, 27132, 26710, 25716, 24288, 22948, 22386, 22256, 22545, 
    22887, 23638, 24658, 25487, 26649, 27216, 27003, 26250, 25778, 25216, 
    24557, 23971,
  27236, 27221, 26956, 26623, 25760, 24359, 22982, 22466, 22313, 22551, 
    22937, 23705, 24628, 25737, 26690, 26914, 26836, 26292, 25851, 25296, 
    24658, 23959,
  27214, 27232, 26794, 26586, 25757, 24435, 23053, 22496, 22298, 22485, 
    22999, 23679, 24673, 25932, 26964, 26584, 26474, 26051, 25685, 25289, 
    24595, 23998,
  27605, 27581, 26710, 26418, 25637, 24425, 23097, 22458, 22255, 22506, 
    22909, 23523, 24515, 25738, 26823, 26379, 25117, 25123, 25141, 24924, 
    24376, 23924,
  27576, 27521, 26799, 26493, 25742, 24512, 23138, 22543, 22273, 22560, 
    22879, 23594, 24574, 25851, 26535, 26489, 25440, 25396, 25216, 24918, 
    24433, 23871,
  27129, 27110, 26912, 26697, 25960, 24637, 23249, 22674, 22332, 22566, 
    22922, 23602, 24511, 25717, 26768, 26660, 26117, 25724, 25463, 25003, 
    24462, 23990,
  27074, 27061, 26980, 26794, 26025, 24779, 23321, 22667, 22418, 22583, 
    22912, 23562, 24480, 25695, 26865, 26952, 26752, 26059, 25632, 25053, 
    24488, 23924,
  26977, 27012, 26988, 26781, 26088, 24789, 23354, 22749, 22426, 22500, 
    22904, 23619, 24504, 25810, 26663, 27188, 27144, 26250, 25609, 25054, 
    24417, 23851,
  26850, 26932, 26897, 26797, 26115, 24848, 23387, 22763, 22395, 22520, 
    22898, 23479, 24562, 25481, 26844, 27213, 27013, 26134, 25572, 24959, 
    24365, 23876,
  26726, 26844, 26839, 26747, 26063, 24853, 23460, 22814, 22458, 22614, 
    22851, 23564, 24445, 25759, 26838, 27151, 26904, 26065, 25570, 25018, 
    24478, 23935,
  26631, 26778, 26816, 26691, 26111, 24885, 23476, 22826, 22469, 22611, 
    22837, 23568, 24393, 25583, 26323, 27101, 26941, 26269, 25676, 25077, 
    24482, 23920,
  26608, 26749, 26706, 26627, 26079, 24918, 23556, 22822, 22500, 22618, 
    22946, 23488, 24348, 25743, 26479, 27089, 27187, 26422, 25874, 25323, 
    24639, 24038,
  26657, 26773, 26738, 26651, 26169, 24976, 23586, 22886, 22480, 22523, 
    22887, 23542, 24464, 25684, 26557, 27100, 27378, 26643, 26112, 25414, 
    24566, 24068,
  26746, 26828, 26774, 26694, 26172, 25008, 23605, 22909, 22505, 22592, 
    22923, 23512, 24342, 25631, 26374, 27105, 27290, 26635, 26088, 25448, 
    24673, 23958,
  26806, 26883, 26779, 26726, 26139, 25042, 23630, 22889, 22501, 22557, 
    22797, 23518, 24368, 25610, 26625, 27040, 26990, 26550, 26088, 25471, 
    24708, 24017,
  26799, 26896, 26685, 26660, 26125, 25062, 23676, 22978, 22536, 22586, 
    22839, 23435, 24448, 25510, 26535, 26920, 27014, 26541, 26026, 25490, 
    24631, 24068,
  26700, 26820, 26640, 26585, 26115, 25037, 23689, 22972, 22596, 22589, 
    22870, 23450, 24442, 25649, 26676, 26795, 26799, 26410, 26026, 25520, 
    24802, 24126,
  26519, 26626, 26469, 26507, 26138, 25061, 23689, 23026, 22540, 22576, 
    22895, 23455, 24271, 25552, 26628, 26717, 26418, 26268, 26006, 25531, 
    24776, 24128,
  26284, 26361, 26451, 26494, 26080, 25104, 23751, 23046, 22666, 22595, 
    22906, 23439, 24390, 25483, 26707, 26722, 26700, 26448, 26110, 25619, 
    24942, 24201,
  26062, 26111, 26376, 26425, 26128, 25119, 23783, 23061, 22624, 22605, 
    22898, 23405, 24239, 25270, 26422, 26788, 26763, 26476, 26075, 25596, 
    24985, 24221,
  25915, 25961, 26334, 26362, 26142, 25145, 23786, 23068, 22649, 22605, 
    22970, 23495, 24348, 25424, 26464, 26789, 26916, 26476, 26147, 25675, 
    24954, 24279,
  25862, 25939, 26279, 26427, 26144, 25161, 23829, 23117, 22646, 22654, 
    22901, 23439, 24362, 25560, 26247, 26825, 26962, 26588, 26225, 25699, 
    24978, 24359,
  25877, 25986, 26320, 26420, 26150, 25181, 23834, 23106, 22704, 22637, 
    22909, 23441, 24315, 25386, 26567, 26804, 27055, 26657, 26334, 25841, 
    25161, 24458,
  25905, 26017, 26328, 26451, 26134, 25179, 23863, 23175, 22692, 22602, 
    22881, 23462, 24428, 25621, 26719, 26750, 27158, 26740, 26360, 25914, 
    25178, 24576,
  25905, 25970, 26317, 26450, 26132, 25194, 23909, 23171, 22683, 22648, 
    22860, 23399, 24281, 25325, 26631, 26578, 26524, 26401, 26150, 25793, 
    25132, 24655,
  25858, 25861, 26318, 26420, 26108, 25245, 23936, 23190, 22753, 22670, 
    22906, 23437, 24325, 25530, 26541, 26613, 26860, 26509, 26224, 25773, 
    25214, 24574,
  25779, 25740, 26246, 26360, 26124, 25231, 23909, 23187, 22712, 22627, 
    22896, 23440, 24317, 25490, 26526, 26674, 27360, 26843, 26406, 25921, 
    25289, 24769,
  25705, 25665, 26199, 26337, 26113, 25276, 23894, 23216, 22725, 22633, 
    22902, 23321, 24168, 25491, 26777, 26691, 27319, 26760, 26349, 25939, 
    25353, 24822,
  25688, 25675, 26099, 26266, 26124, 25224, 23888, 23181, 22749, 22661, 
    22934, 23345, 24132, 25335, 26840, 26579, 27175, 26726, 26359, 25937, 
    25493, 24898,
  25784, 25819, 26134, 26244, 26089, 25212, 23928, 23203, 22790, 22626, 
    22844, 23475, 24177, 25326, 26425, 26487, 27131, 26666, 26281, 25950, 
    25550, 25153,
  26008, 26100, 26237, 26338, 26019, 25200, 23912, 23193, 22786, 22687, 
    22988, 23483, 24274, 25414, 26307, 26576, 26896, 26497, 26240, 25918, 
    25525, 25159,
  26320, 26457, 26464, 26510, 26132, 25264, 23971, 23212, 22828, 22712, 
    22857, 23476, 24201, 25419, 26191, 26704, 26809, 26395, 26100, 25782, 
    25429, 25031,
  26625, 26792, 26640, 26528, 26144, 25182, 23959, 23243, 22835, 22676, 
    22888, 23357, 24155, 25501, 26651, 26743, 26760, 26356, 26066, 25745, 
    25428, 24937,
  26833, 27027, 26617, 26591, 26163, 25226, 23953, 23245, 22793, 22726, 
    22938, 23407, 24178, 25406, 26550, 26746, 26694, 26253, 25954, 25566, 
    25256, 24964,
  26920, 27155, 26716, 26613, 26194, 25250, 23945, 23298, 22876, 22688, 
    22910, 23358, 24142, 25437, 26765, 26683, 26044, 25718, 25486, 25259, 
    24880, 24510,
  26935, 27199, 26697, 26586, 26166, 25272, 23980, 23298, 22830, 22745, 
    22904, 23455, 24223, 25404, 26391, 26734, 26085, 25644, 25382, 25091, 
    24720, 24403,
  26931, 27201, 26642, 26639, 26210, 25277, 24001, 23308, 22856, 22644, 
    22882, 23382, 24372, 25257, 26596, 26718, 26641, 25994, 25638, 25246, 
    24828, 24398,
  26927, 27168, 26677, 26599, 26198, 25311, 24004, 23297, 22894, 22737, 
    22937, 23372, 24190, 25312, 26729, 26675, 26485, 25982, 25672, 25352, 
    24880, 24521,
  26889, 27082, 26575, 26585, 26189, 25285, 24006, 23295, 22879, 22737, 
    23027, 23396, 24308, 25510, 26876, 26632, 25972, 25656, 25347, 25183, 
    24765, 24374,
  26768, 26918, 26616, 26613, 26213, 25293, 24015, 23326, 22899, 22726, 
    22911, 23287, 24258, 25453, 26056, 26621, 25963, 25526, 25283, 24978, 
    24717, 24268,
  26531, 26672, 26600, 26554, 26206, 25311, 24010, 23303, 22841, 22691, 
    22989, 23339, 24075, 25416, 26481, 26635, 26732, 26069, 25725, 25266, 
    24837, 24323,
  26177, 26332, 26425, 26565, 26203, 25306, 24009, 23340, 22898, 22723, 
    22931, 23457, 24229, 25260, 26856, 26660, 26765, 26175, 25755, 25341, 
    24781, 24476,
  25710, 25899, 26312, 26432, 26179, 25327, 24034, 23359, 22886, 22784, 
    23032, 23447, 24260, 25334, 26859, 26482, 26785, 26204, 25712, 25254, 
    24761, 24416,
  25196, 25410, 26022, 26276, 26109, 25261, 24006, 23311, 22925, 22732, 
    22925, 23423, 24275, 25319, 26510, 26167, 26637, 26123, 25668, 25292, 
    24704, 24315,
  24726, 24950, 25723, 26069, 25985, 25240, 24056, 23378, 22925, 22757, 
    22962, 23306, 24312, 25314, 26532, 25840, 26493, 26317, 25755, 25282, 
    24736, 24327,
  24425, 24631, 25591, 26021, 26027, 25256, 24043, 23324, 22929, 22810, 
    22975, 23421, 24256, 25158, 26476, 25673, 26863, 26542, 26013, 25382, 
    24849, 24279,
  24345, 24530, 25584, 26021, 26003, 25301, 24009, 23391, 22887, 22744, 
    22975, 23451, 24163, 25317, 26739, 25646, 26997, 26822, 26231, 25609, 
    24925, 24425,
  24460, 24642, 25797, 26128, 26052, 25295, 24040, 23333, 22925, 22714, 
    22895, 23487, 24292, 25411, 26474, 25819, 27226, 26913, 26284, 25769, 
    25008, 24517,
  24654, 24865, 26021, 26225, 26149, 25290, 23991, 23320, 22899, 22765, 
    22917, 23401, 24201, 25287, 26461, 26159, 27301, 26929, 26356, 25751, 
    25097, 24504,
  24817, 25054, 26125, 26301, 26103, 25307, 24031, 23361, 22898, 22809, 
    22979, 23507, 24215, 25324, 26644, 26312, 27344, 26903, 26353, 25735, 
    25057, 24478,
  24847, 25087, 26209, 26359, 26165, 25259, 24002, 23323, 22937, 22811, 
    22958, 23345, 24333, 25549, 26379, 26459, 27357, 26904, 26384, 25813, 
    25103, 24498,
  24681, 24903, 26229, 26371, 26141, 25289, 24007, 23371, 22940, 22821, 
    22981, 23388, 24276, 25476, 26531, 26551, 27459, 26972, 26401, 25797, 
    25071, 24465,
  24305, 24531, 26078, 26197, 26114, 25293, 23987, 23297, 22919, 22809, 
    22967, 23466, 24299, 25593, 26779, 26351, 27453, 26891, 26408, 25828, 
    25109, 24460,
  23731, 24005, 25666, 25976, 25908, 25183, 23976, 23362, 22945, 22744, 
    22988, 23492, 24171, 25282, 26538, 26015, 27266, 26940, 26363, 25878, 
    25148, 24479,
  22999, 23346, 25207, 25604, 25801, 25151, 23970, 23328, 22959, 22771, 
    22897, 23408, 24218, 25331, 26901, 25628, 27091, 26887, 26368, 25868, 
    25256, 24540,
  22196, 22592, 24670, 25262, 25613, 25113, 23960, 23349, 22914, 22883, 
    22970, 23406, 24321, 25382, 26360, 24984, 26720, 26813, 26362, 25918, 
    25155, 24594,
  21436, 21865, 23862, 24794, 25372, 25019, 23958, 23376, 22937, 22808, 
    23007, 23462, 24314, 25427, 26661, 24035, 26026, 26710, 26334, 25898, 
    25137, 24628,
  20851, 21284, 23559, 24529, 25292, 25025, 23915, 23347, 22947, 22807, 
    23023, 23407, 24246, 25496, 26574, 23436, 25784, 26707, 26401, 25987, 
    25310, 24581,
  20562, 20967, 23668, 24646, 25336, 25028, 23933, 23312, 22939, 22821, 
    22992, 23514, 24280, 25275, 26596, 23490, 25954, 26682, 26434, 25985, 
    25254, 24689,
  20592, 20967, 23893, 24765, 25337, 24978, 23940, 23318, 22983, 22832, 
    23061, 23362, 24302, 25377, 26551, 23804, 26101, 26724, 26428, 25937, 
    25255, 24737,
  20885, 21245, 23966, 24778, 25348, 24965, 23878, 23290, 22950, 22818, 
    23061, 23492, 24204, 25370, 26963, 23909, 26163, 26685, 26353, 25969, 
    25263, 24667,
  21330, 21661, 23988, 24821, 25341, 24976, 23878, 23285, 22968, 22852, 
    23001, 23512, 24314, 25399, 26472, 23893, 25814, 26662, 26367, 25951, 
    25334, 24776,
  21772, 22052, 24206, 24926, 25395, 24928, 23886, 23280, 22933, 22839, 
    23064, 23461, 24210, 25430, 26817, 24043, 25927, 26734, 26395, 25938, 
    25264, 24764,
  22084, 22316, 24303, 24980, 25408, 24897, 23876, 23251, 22943, 22827, 
    22987, 23490, 24276, 25528, 26668, 24129, 25876, 26712, 26357, 25900, 
    25276, 24710,
  22229, 22445, 24287, 25002, 25383, 24909, 23837, 23295, 22998, 22923, 
    23066, 23453, 24287, 25495, 26661, 24048, 25868, 26595, 26304, 25899, 
    25253, 24743,
  22234, 22458, 24204, 24961, 25379, 24910, 23854, 23249, 22990, 22878, 
    23032, 23493, 24350, 25475, 27089, 23954, 25850, 26598, 26332, 25839, 
    25215, 24679,
  22134, 22354, 24120, 24936, 25394, 24891, 23847, 23309, 22995, 22872, 
    22989, 23460, 24354, 25610, 26660, 23910, 25940, 26556, 26331, 25850, 
    25242, 24727,
  21921, 22118, 24147, 25003, 25422, 24876, 23801, 23266, 22953, 22926, 
    23061, 23466, 24443, 25665, 26621, 24178, 26138, 26647, 26335, 25791, 
    25218, 24802,
  21568, 21763, 24013, 24888, 25360, 24816, 23774, 23282, 23015, 22905, 
    22995, 23549, 24312, 25554, 26956, 24131, 26061, 26563, 26316, 25836, 
    25208, 24830,
  21127, 21352, 23617, 24656, 25264, 24807, 23747, 23278, 22958, 22876, 
    23127, 23558, 24455, 25451, 26602, 23710, 25884, 26606, 26262, 25840, 
    25284, 24761,
  20742, 21013, 23372, 24569, 25178, 24728, 23718, 23240, 23015, 22911, 
    23103, 23468, 24374, 25480, 26711, 23362, 25763, 26453, 26170, 25747, 
    25293, 24676,
  20588, 20874, 23459, 24548, 25199, 24726, 23735, 23228, 22987, 22910, 
    23067, 23531, 24451, 25679, 26773, 23469, 25885, 26464, 26087, 25596, 
    25097, 24669,
  20726, 21005, 23684, 24693, 25212, 24777, 23745, 23271, 22990, 22917, 
    23087, 23570, 24284, 25549, 26625, 23746, 25977, 26440, 26066, 25661, 
    25073, 24610,
  21072, 21337, 23890, 24850, 25287, 24744, 23710, 23256, 23057, 22951, 
    23122, 23654, 24512, 25873, 27023, 24099, 26083, 26525, 26184, 25704, 
    25093, 24485,
  21423, 21725, 24162, 24945, 25321, 24670, 23679, 23227, 23037, 22939, 
    23130, 23712, 24427, 25819, 26954, 24361, 26184, 26472, 26122, 25664, 
    25113, 24611,
  21646, 22004, 24303, 25059, 25309, 24684, 23653, 23234, 23035, 22940, 
    23211, 23572, 24442, 25640, 27153, 24461, 26278, 26534, 26161, 25735, 
    25089, 24525,
  21699, 22107, 24422, 25098, 25318, 24622, 23687, 23251, 23043, 22970, 
    23251, 23701, 24413, 25772, 26965, 24514, 26284, 26444, 26163, 25687, 
    25034, 24493,
  21685, 22068, 24443, 25103, 25298, 24628, 23643, 23234, 23016, 22979, 
    23128, 23632, 24435, 25674, 26963, 24422, 26200, 26476, 26123, 25670, 
    25137, 24615,
  21678, 22023, 24449, 25141, 25307, 24593, 23597, 23251, 22985, 23003, 
    23113, 23640, 24440, 25769, 26959, 24326, 26115, 26481, 26077, 25740, 
    25102, 24529,
  21747, 22043, 24435, 25129, 25273, 24563, 23564, 23229, 23069, 22989, 
    23199, 23706, 24528, 25910, 26919, 24186, 26091, 26462, 26197, 25830, 
    25300, 24584,
  21882, 22140, 24430, 25142, 25271, 24550, 23576, 23203, 23079, 22992, 
    23117, 23663, 24505, 26029, 26926, 24149, 26000, 26457, 26150, 25794, 
    25268, 24592,
  22057, 22276, 24486, 25144, 25251, 24483, 23543, 23241, 23076, 23007, 
    23260, 23607, 24684, 25813, 26834, 24096, 26004, 26456, 26171, 25830, 
    25224, 24726,
  22234, 22436, 24570, 25187, 25260, 24462, 23537, 23213, 23027, 23027, 
    23161, 23633, 24665, 25778, 26891, 24134, 26035, 26395, 26103, 25762, 
    25167, 24715,
  22429, 22613, 24645, 25264, 25273, 24434, 23525, 23201, 23105, 23087, 
    23083, 23740, 24715, 25609, 26688, 24254, 26199, 26475, 26115, 25719, 
    25104, 24468,
  22648, 22817, 24843, 25372, 25243, 24422, 23531, 23195, 23127, 23073, 
    23218, 23657, 24656, 25832, 27079, 24372, 26226, 26388, 26086, 25648, 
    25060, 24583,
  22904, 23052, 24989, 25441, 25260, 24393, 23511, 23212, 23090, 23103, 
    23227, 23693, 24628, 25843, 26772, 24493, 26359, 26360, 26029, 25753, 
    25169, 24563,
  23192, 23312, 25161, 25530, 25161, 24334, 23474, 23213, 23082, 23043, 
    23244, 23787, 24747, 25823, 26950, 24664, 26332, 26298, 26025, 25654, 
    25125, 24469,
  23493, 23583, 25301, 25535, 25186, 24299, 23428, 23212, 23101, 23063, 
    23282, 23821, 24721, 26059, 27531, 24669, 26234, 26303, 25963, 25575, 
    25011, 24416,
  23785, 23829, 25399, 25533, 25122, 24230, 23402, 23200, 23160, 23095, 
    23288, 23824, 24826, 26029, 27053, 24550, 26169, 26208, 25824, 25448, 
    24925, 24297,
  24037, 24037, 25411, 25542, 25070, 24159, 23380, 23216, 23142, 23074, 
    23335, 23877, 24739, 26096, 26979, 24483, 26132, 26188, 25737, 25384, 
    24812, 24233,
  24136, 24105, 25509, 25554, 25032, 24147, 23350, 23188, 23114, 23041, 
    23357, 23883, 25010, 26143, 27271, 24590, 26063, 26095, 25770, 25343, 
    24776, 24249,
  23997, 23948, 25525, 25576, 25008, 24067, 23354, 23201, 23161, 23148, 
    23310, 23883, 24856, 26272, 27083, 24718, 26183, 26035, 25688, 25253, 
    24741, 24146,
  23651, 23613, 25614, 25529, 24912, 23985, 23326, 23211, 23144, 23103, 
    23284, 23870, 24893, 26038, 27200, 24866, 26268, 25971, 25560, 25125, 
    24603, 24035,
  23477, 23430, 25565, 25500, 24873, 23925, 23300, 23150, 23076, 23072, 
    23282, 23955, 25048, 26311, 27015, 24910, 26363, 25932, 25512, 25045, 
    24432, 23943,
  27331, 27305, 27308, 26835, 25695, 24114, 22762, 22345, 22278, 22559, 
    22939, 23709, 24765, 26010, 26911, 27696, 27104, 26172, 25524, 25037, 
    24253, 23714,
  27309, 27277, 27329, 26844, 25763, 24261, 22895, 22389, 22298, 22570, 
    22917, 23686, 24685, 25815, 26701, 27584, 27163, 26148, 25572, 24976, 
    24379, 23794,
  27265, 27235, 27069, 26681, 25688, 24305, 22926, 22412, 22275, 22495, 
    22974, 23680, 24573, 25776, 26759, 27211, 26950, 26186, 25685, 25076, 
    24413, 23701,
  27203, 27196, 26838, 26553, 25703, 24365, 23005, 22454, 22322, 22513, 
    22981, 23587, 24515, 25963, 26553, 26766, 26621, 26177, 25694, 25162, 
    24502, 23875,
  27203, 27216, 26757, 26493, 25686, 24374, 23080, 22482, 22319, 22590, 
    23024, 23570, 24526, 25619, 26725, 26406, 25848, 25670, 25399, 24962, 
    24337, 23672,
  27615, 27579, 26714, 26367, 25651, 24445, 23089, 22493, 22227, 22459, 
    22870, 23522, 24496, 25578, 26266, 26478, 24989, 25101, 25060, 24840, 
    24214, 23820,
  27185, 27200, 26888, 26681, 25913, 24529, 23167, 22588, 22351, 22559, 
    22926, 23553, 24425, 25668, 26769, 26716, 26388, 25863, 25474, 25013, 
    24439, 23773,
  27148, 27166, 27026, 26814, 26032, 24659, 23265, 22626, 22359, 22545, 
    22923, 23571, 24494, 25722, 26939, 27120, 27078, 26163, 25589, 24994, 
    24356, 23725,
  27095, 27147, 27036, 26882, 26074, 24751, 23289, 22726, 22399, 22585, 
    22903, 23493, 24601, 25705, 26588, 27302, 27165, 26182, 25524, 24975, 
    24306, 23692,
  27012, 27111, 27078, 26860, 26144, 24767, 23360, 22714, 22418, 22559, 
    22874, 23461, 24414, 25632, 26395, 27369, 27159, 26121, 25542, 24938, 
    24274, 23653,
  26903, 27031, 26982, 26830, 26147, 24823, 23411, 22787, 22449, 22590, 
    22901, 23537, 24461, 25786, 26966, 27324, 27022, 25975, 25415, 24837, 
    24279, 23737,
  26783, 26933, 26916, 26751, 26116, 24859, 23439, 22773, 22441, 22570, 
    22972, 23550, 24472, 25764, 26565, 27266, 26957, 26138, 25510, 24927, 
    24290, 23763,
  26668, 26848, 26815, 26704, 26072, 24896, 23461, 22826, 22494, 22569, 
    22887, 23553, 24442, 25615, 26858, 27138, 27056, 26335, 25775, 25104, 
    24415, 23909,
  26609, 26787, 26685, 26693, 26157, 24961, 23517, 22863, 22478, 22540, 
    22933, 23586, 24456, 25495, 26601, 27165, 27283, 26531, 25937, 25282, 
    24489, 23947,
  26623, 26770, 26726, 26646, 26156, 25007, 23536, 22880, 22541, 22562, 
    22880, 23472, 24334, 25543, 26488, 27141, 27374, 26725, 26169, 25435, 
    24581, 23903,
  26689, 26795, 26760, 26657, 26113, 24949, 23601, 22920, 22515, 22542, 
    22916, 23412, 24439, 25663, 26586, 27111, 27236, 26644, 26146, 25501, 
    24593, 23880,
  26745, 26840, 26715, 26679, 26123, 24986, 23636, 22907, 22543, 22536, 
    22892, 23444, 24410, 25425, 26743, 27027, 27123, 26529, 26056, 25400, 
    24622, 23918,
  26753, 26851, 26753, 26653, 26121, 25034, 23678, 22945, 22581, 22594, 
    22894, 23434, 24468, 25557, 26750, 26973, 27117, 26484, 26021, 25393, 
    24589, 23970,
  26678, 26777, 26577, 26626, 26113, 25022, 23674, 22957, 22598, 22585, 
    22883, 23559, 24362, 25545, 26688, 26882, 27045, 26513, 26124, 25504, 
    24798, 23976,
  26523, 26598, 26496, 26553, 26113, 25055, 23695, 22979, 22594, 22565, 
    22797, 23434, 24380, 25706, 26699, 26804, 26919, 26507, 26124, 25584, 
    24862, 24205,
  26312, 26370, 26409, 26479, 26118, 25096, 23692, 23031, 22614, 22611, 
    22890, 23404, 24232, 25600, 26783, 26793, 27039, 26615, 26168, 25660, 
    24951, 24271,
  26121, 26179, 26390, 26416, 26091, 25116, 23743, 23037, 22631, 22621, 
    22987, 23460, 24451, 25382, 26431, 26834, 27116, 26641, 26215, 25704, 
    25065, 24244,
  26016, 26084, 26348, 26423, 26151, 25171, 23778, 23035, 22637, 22632, 
    22843, 23506, 24415, 25629, 27034, 26815, 27050, 26665, 26162, 25716, 
    25040, 24236,
  26003, 26097, 26294, 26441, 26139, 25127, 23801, 23082, 22682, 22679, 
    22965, 23355, 24307, 25424, 26638, 26823, 27071, 26581, 26232, 25744, 
    25127, 24442,
  26048, 26158, 26385, 26459, 26136, 25162, 23815, 23121, 22672, 22582, 
    22879, 23455, 24227, 25266, 26444, 26773, 27213, 26693, 26322, 25800, 
    25093, 24494,
  26087, 26192, 26365, 26478, 26151, 25185, 23890, 23117, 22708, 22635, 
    22885, 23471, 24286, 25375, 26525, 26734, 26998, 26560, 26238, 25768, 
    25161, 24445,
  26073, 26141, 26311, 26440, 26166, 25172, 23828, 23174, 22725, 22650, 
    22842, 23336, 24289, 25545, 26664, 26688, 26864, 26496, 26138, 25690, 
    25090, 24457,
  25993, 26017, 26281, 26394, 26091, 25203, 23921, 23149, 22733, 22692, 
    22899, 23367, 24323, 25303, 26378, 26724, 27293, 26719, 26238, 25819, 
    25261, 24705,
  25868, 25864, 26178, 26385, 26090, 25178, 23853, 23202, 22712, 22681, 
    22897, 23427, 24290, 25604, 26539, 26646, 27307, 26691, 26284, 25868, 
    25336, 24792,
  25741, 25740, 25990, 26235, 26063, 25201, 23893, 23172, 22762, 22703, 
    22869, 23400, 24258, 25263, 26590, 26499, 27191, 26653, 26337, 25861, 
    25406, 24899,
  25667, 25692, 25901, 26168, 26053, 25204, 23898, 23236, 22811, 22672, 
    22961, 23404, 24192, 25277, 26971, 26379, 27097, 26649, 26244, 25846, 
    25450, 24981,
  25713, 25777, 25993, 26197, 26030, 25181, 23947, 23218, 22773, 22694, 
    22880, 23403, 24198, 25141, 26614, 26429, 26960, 26472, 26159, 25803, 
    25394, 25108,
  25914, 26016, 26206, 26318, 26037, 25169, 23914, 23196, 22769, 22660, 
    22879, 23373, 24249, 25268, 26546, 26510, 26886, 26425, 26083, 25715, 
    25432, 24961,
  26243, 26363, 26498, 26432, 26116, 25203, 23911, 23193, 22785, 22665, 
    22895, 23339, 24299, 25271, 26454, 26716, 26968, 26381, 26040, 25617, 
    25203, 24934,
  26604, 26734, 26646, 26567, 26148, 25216, 23944, 23210, 22812, 22629, 
    22830, 23379, 24296, 25160, 26402, 26826, 26944, 26385, 25950, 25604, 
    25157, 24779,
  26884, 27038, 26671, 26600, 26199, 25192, 23966, 23260, 22835, 22644, 
    22931, 23375, 24109, 25206, 26546, 26838, 26926, 26312, 25874, 25488, 
    25004, 24538,
  27035, 27240, 26724, 26605, 26218, 25225, 23979, 23238, 22819, 22690, 
    23037, 23395, 24195, 25150, 26732, 26793, 26520, 26137, 25825, 25380, 
    24978, 24520,
  27082, 27330, 26734, 26605, 26185, 25247, 23965, 23281, 22766, 22727, 
    22993, 23284, 24265, 25334, 26201, 26771, 26750, 26200, 25763, 25337, 
    24901, 24560,
  27067, 27330, 26734, 26599, 26212, 25258, 23990, 23258, 22831, 22735, 
    22955, 23435, 24175, 25693, 26592, 26810, 26881, 26291, 25825, 25336, 
    24888, 24522,
  27005, 27239, 26684, 26565, 26207, 25224, 23985, 23300, 22854, 22639, 
    22882, 23422, 24195, 25362, 26375, 26734, 26756, 26250, 25784, 25411, 
    24902, 24443,
  26860, 27039, 26747, 26601, 26233, 25265, 23998, 23301, 22856, 22667, 
    22960, 23396, 24331, 25434, 26657, 26739, 26624, 26018, 25693, 25242, 
    24787, 24410,
  26583, 26706, 26615, 26608, 26245, 25237, 23987, 23317, 22888, 22704, 
    22879, 23440, 24243, 25419, 26429, 26722, 27019, 26263, 25789, 25280, 
    24796, 24231,
  26150, 26250, 26438, 26501, 26201, 25258, 24051, 23303, 22845, 22733, 
    22962, 23376, 24324, 25454, 26482, 26691, 26735, 26028, 25595, 25138, 
    24655, 24251,
  25591, 25698, 26160, 26340, 26123, 25311, 23960, 23260, 22899, 22736, 
    22895, 23383, 24333, 25442, 26313, 26372, 26532, 25988, 25598, 25188, 
    24726, 24204,
  24964, 25099, 25744, 26099, 26019, 25271, 24001, 23338, 22872, 22780, 
    22970, 23412, 24203, 25354, 26527, 25967, 26682, 26212, 25748, 25232, 
    24706, 24137,
  24372, 24535, 25460, 25878, 25941, 25241, 24022, 23313, 22905, 22691, 
    22951, 23405, 24164, 25280, 26324, 25632, 26657, 26363, 25869, 25307, 
    24866, 24292,
  23910, 24094, 25272, 25751, 25903, 25198, 24031, 23309, 22905, 22750, 
    22845, 23369, 24041, 25421, 26639, 25333, 26726, 26548, 26061, 25458, 
    24936, 24397,
  23664, 23844, 25130, 25734, 25933, 25237, 24001, 23332, 22888, 22726, 
    22933, 23405, 24304, 25452, 26500, 25180, 26717, 26818, 26257, 25634, 
    24947, 24335,
  23637, 23801, 25296, 25822, 25935, 25240, 24018, 23302, 22864, 22776, 
    22953, 23359, 24203, 25490, 26638, 25379, 26963, 26888, 26432, 25749, 
    25074, 24528,
  23754, 23909, 25570, 25987, 25978, 25261, 24014, 23300, 22937, 22747, 
    22979, 23379, 24262, 25250, 26290, 25790, 27291, 26907, 26342, 25797, 
    25151, 24567,
  23873, 24051, 25760, 26035, 25995, 25290, 23979, 23320, 22955, 22745, 
    22965, 23410, 24197, 25287, 26683, 26006, 27417, 26938, 26420, 25872, 
    25093, 24527,
  23895, 24101, 25718, 26070, 26015, 25248, 23999, 23320, 22904, 22782, 
    22998, 23460, 24346, 25408, 26326, 26112, 27347, 27026, 26391, 25769, 
    25047, 24468,
  23760, 23983, 25657, 25979, 25975, 25259, 23970, 23296, 22854, 22790, 
    22936, 23326, 24344, 25429, 26604, 26059, 27279, 26964, 26393, 25828, 
    25131, 24568,
  23459, 23679, 25535, 25957, 25907, 25208, 23982, 23297, 22940, 22740, 
    22995, 23224, 24308, 25285, 26637, 26037, 27350, 26944, 26417, 25893, 
    25106, 24568,
  23019, 23255, 25143, 25648, 25783, 25147, 23955, 23279, 22905, 22785, 
    22969, 23412, 24174, 25314, 26773, 25680, 27363, 27016, 26451, 25893, 
    25170, 24589,
  22488, 22772, 24604, 25304, 25637, 25126, 23961, 23298, 22935, 22769, 
    22936, 23412, 24278, 25434, 26885, 25008, 26759, 26847, 26421, 25868, 
    25176, 24542,
  21932, 22271, 24249, 24993, 25476, 25045, 23931, 23315, 22942, 22813, 
    22984, 23425, 24174, 25406, 26641, 24540, 26434, 26722, 26363, 25832, 
    25240, 24495,
  21427, 21789, 23915, 24821, 25373, 24989, 23935, 23301, 22920, 22819, 
    23022, 23369, 24211, 25312, 26597, 24118, 26075, 26670, 26335, 25776, 
    25100, 24443,
  21041, 21409, 23657, 24640, 25289, 24952, 23913, 23335, 22976, 22787, 
    22911, 23383, 24268, 25488, 26470, 23642, 26029, 26711, 26350, 25932, 
    25184, 24624,
  20825, 21182, 23545, 24605, 25262, 24929, 23921, 23291, 22936, 22855, 
    23024, 23485, 24251, 25254, 26636, 23453, 25924, 26737, 26403, 25953, 
    25274, 24711,
  20821, 21152, 23740, 24674, 25273, 24907, 23883, 23286, 22960, 22803, 
    23090, 23439, 24339, 25236, 26569, 23666, 25957, 26728, 26415, 26025, 
    25314, 24692,
  21005, 21322, 23911, 24765, 25315, 24962, 23898, 23250, 22948, 22848, 
    23006, 23493, 24423, 25224, 26610, 23957, 26116, 26725, 26429, 26071, 
    25297, 24713,
  21317, 21644, 23899, 24784, 25337, 24951, 23836, 23273, 22945, 22823, 
    22979, 23368, 24306, 25387, 26572, 23923, 25979, 26629, 26403, 25941, 
    25253, 24711,
  21691, 22008, 23879, 24832, 25327, 24922, 23857, 23293, 22978, 22914, 
    22965, 23410, 24322, 25346, 26889, 23810, 25873, 26699, 26424, 26004, 
    25368, 24773,
  22039, 22317, 24210, 24982, 25382, 24945, 23875, 23262, 22966, 22870, 
    23074, 23453, 24284, 25375, 26417, 24041, 25961, 26691, 26431, 25991, 
    25362, 24807,
  22288, 22521, 24367, 25096, 25422, 24914, 23858, 23299, 22976, 22858, 
    23017, 23385, 24338, 25478, 26659, 24175, 26015, 26625, 26352, 25891, 
    25293, 24740,
  22408, 22627, 24417, 25087, 25399, 24839, 23832, 23283, 22963, 22845, 
    23068, 23569, 24349, 25163, 26601, 24178, 25957, 26654, 26313, 25946, 
    25262, 24712,
  22401, 22634, 24281, 25013, 25392, 24882, 23797, 23270, 22962, 22876, 
    23042, 23561, 24387, 25415, 26864, 24128, 26100, 26635, 26300, 25768, 
    25237, 24682,
  22274, 22511, 24202, 25033, 25386, 24815, 23774, 23253, 22978, 22932, 
    23113, 23505, 24291, 25440, 26600, 24154, 26103, 26579, 26340, 25802, 
    25296, 24777,
  22015, 22227, 24280, 25012, 25342, 24826, 23776, 23257, 22968, 22978, 
    22985, 23511, 24367, 25421, 26954, 24301, 26178, 26625, 26324, 25843, 
    25354, 24785,
  21606, 21805, 24021, 24886, 25320, 24814, 23807, 23255, 22993, 22956, 
    23082, 23584, 24468, 25491, 26607, 24123, 26138, 26651, 26228, 25801, 
    25306, 24786,
  21122, 21345, 23767, 24692, 25224, 24774, 23778, 23249, 22990, 22943, 
    23111, 23509, 24293, 25591, 26671, 23810, 26005, 26600, 26236, 25718, 
    25230, 24696,
  20720, 20997, 23555, 24603, 25264, 24759, 23769, 23256, 23007, 22922, 
    23070, 23604, 24360, 25538, 26756, 23604, 25847, 26540, 26131, 25626, 
    25181, 24632,
  20579, 20890, 23526, 24581, 25168, 24740, 23741, 23245, 23014, 23015, 
    23145, 23574, 24460, 25532, 27022, 23617, 25957, 26458, 26013, 25581, 
    25074, 24478,
  20748, 21067, 23643, 24618, 25175, 24701, 23687, 23256, 23001, 22950, 
    23063, 23561, 24523, 25427, 26532, 23791, 26018, 26434, 26068, 25607, 
    24962, 24519,
  21143, 21438, 23861, 24757, 25239, 24676, 23695, 23226, 23005, 22942, 
    23084, 23626, 24478, 25490, 26944, 24049, 26086, 26489, 26130, 25621, 
    25070, 24655,
  21561, 21863, 24069, 24905, 25243, 24676, 23657, 23232, 22965, 23032, 
    23112, 23622, 24380, 25492, 26781, 24255, 26093, 26466, 26172, 25748, 
    25148, 24567,
  21863, 22190, 24269, 25036, 25258, 24673, 23655, 23204, 23054, 23031, 
    23212, 23696, 24423, 25697, 26899, 24450, 26119, 26434, 26135, 25626, 
    25060, 24548,
  21990, 22351, 24400, 25072, 25304, 24640, 23669, 23230, 23023, 22954, 
    23171, 23695, 24544, 25648, 26886, 24543, 26231, 26453, 26151, 25603, 
    24961, 24576,
  22017, 22362, 24412, 25050, 25292, 24609, 23670, 23195, 23055, 22976, 
    23178, 23639, 24440, 25744, 26699, 24433, 26203, 26512, 26214, 25673, 
    25153, 24537,
  22009, 22341, 24392, 25086, 25291, 24591, 23623, 23239, 23041, 22945, 
    23145, 23723, 24365, 25709, 26996, 24312, 26049, 26497, 26183, 25731, 
    25219, 24712,
  22034, 22345, 24413, 25117, 25251, 24586, 23591, 23196, 23043, 23083, 
    23112, 23809, 24521, 25557, 26890, 24287, 26050, 26515, 26212, 25839, 
    25303, 24607,
  22092, 22385, 24441, 25186, 25266, 24506, 23596, 23200, 23047, 23071, 
    23178, 23667, 24577, 25912, 26901, 24270, 26096, 26451, 26200, 25828, 
    25207, 24688,
  22173, 22433, 24495, 25169, 25231, 24458, 23542, 23194, 23079, 23083, 
    23198, 23746, 24524, 25743, 26816, 24207, 26107, 26442, 26207, 25678, 
    25226, 24650,
  22262, 22500, 24594, 25212, 25255, 24460, 23522, 23189, 23045, 23017, 
    23197, 23719, 24607, 25996, 26963, 24246, 26119, 26425, 26166, 25740, 
    25119, 24638,
  22400, 22611, 24707, 25262, 25245, 24409, 23526, 23193, 23126, 23057, 
    23212, 23750, 24609, 25891, 26743, 24371, 26196, 26411, 26048, 25653, 
    25017, 24364,
  22604, 22792, 24887, 25370, 25212, 24392, 23513, 23224, 23081, 23038, 
    23231, 23864, 24553, 25832, 27016, 24514, 26441, 26382, 26095, 25701, 
    25101, 24472,
  22883, 23045, 25041, 25431, 25192, 24348, 23451, 23188, 23088, 23139, 
    23211, 23737, 24629, 26048, 26987, 24689, 26399, 26404, 26073, 25694, 
    25045, 24553,
  23213, 23346, 25154, 25493, 25173, 24264, 23460, 23210, 23074, 23107, 
    23115, 23794, 24659, 25703, 26934, 24801, 26347, 26313, 26041, 25570, 
    25026, 24499,
  23547, 23654, 25312, 25474, 25175, 24246, 23410, 23174, 23155, 23039, 
    23264, 23756, 24817, 26075, 26948, 24811, 26324, 26332, 25932, 25472, 
    24894, 24312,
  23844, 23908, 25314, 25601, 25137, 24194, 23408, 23197, 23094, 23045, 
    23218, 23729, 24612, 26007, 26788, 24567, 26215, 26252, 25895, 25475, 
    24857, 24326,
  24076, 24088, 25369, 25508, 25093, 24142, 23421, 23192, 23143, 23096, 
    23265, 23871, 24720, 26131, 26935, 24421, 26023, 26204, 25863, 25387, 
    24860, 24356,
  24154, 24118, 25323, 25525, 25001, 24094, 23339, 23146, 23156, 23086, 
    23317, 23821, 24937, 26126, 27279, 24417, 26060, 26175, 25758, 25295, 
    24848, 24252,
  24013, 23946, 25415, 25501, 24972, 24042, 23328, 23215, 23098, 23159, 
    23348, 23917, 24857, 26329, 27120, 24481, 26092, 26079, 25690, 25218, 
    24724, 24195,
  23680, 23622, 25445, 25471, 24904, 24010, 23310, 23164, 23151, 23082, 
    23391, 23899, 25043, 26398, 27133, 24604, 26071, 26031, 25665, 25214, 
    24555, 24192,
  23514, 23449, 25498, 25514, 24831, 23903, 23278, 23168, 23121, 23169, 
    23362, 23913, 25027, 26392, 27251, 24765, 26248, 25963, 25542, 25042, 
    24530, 23966,
  27310, 27265, 27328, 26795, 25651, 24150, 22768, 22329, 22254, 22537, 
    22948, 23745, 24690, 25988, 26866, 27635, 27065, 26099, 25551, 24935, 
    24317, 23811,
  27286, 27240, 27261, 26860, 25704, 24232, 22837, 22391, 22242, 22618, 
    22995, 23708, 24668, 25728, 26525, 27610, 27210, 26212, 25656, 25128, 
    24406, 23757,
  27241, 27206, 26986, 26657, 25721, 24313, 22944, 22402, 22234, 22552, 
    22918, 23554, 24567, 25774, 26599, 27250, 27065, 26286, 25685, 25154, 
    24331, 23857,
  27182, 27175, 26843, 26591, 25707, 24372, 23006, 22444, 22293, 22579, 
    22896, 23624, 24525, 25837, 26653, 26788, 26506, 26010, 25591, 25109, 
    24350, 23798,
  27194, 27199, 26747, 26512, 25721, 24429, 23085, 22569, 22307, 22552, 
    23024, 23562, 24567, 25933, 26646, 26593, 26014, 25785, 25454, 24953, 
    24287, 23622,
  27212, 27219, 26941, 26639, 25797, 24505, 23142, 22566, 22340, 22625, 
    22874, 23579, 24600, 25863, 26462, 26760, 26590, 25945, 25496, 24885, 
    24261, 23655,
  27202, 27207, 27065, 26815, 26010, 24571, 23214, 22599, 22410, 22573, 
    22987, 23501, 24572, 25904, 26884, 27129, 27051, 26085, 25460, 24860, 
    24281, 23770,
  27167, 27198, 27138, 26937, 26076, 24667, 23252, 22654, 22388, 22571, 
    22895, 23580, 24593, 25609, 26751, 27335, 27212, 26040, 25465, 24916, 
    24274, 23735,
  27117, 27196, 27109, 26907, 26118, 24708, 23277, 22660, 22390, 22585, 
    22958, 23568, 24448, 25718, 26696, 27410, 26901, 25900, 25379, 24865, 
    24243, 23715,
  27047, 27163, 27057, 26908, 26165, 24801, 23365, 22728, 22446, 22579, 
    22943, 23541, 24544, 25876, 27045, 27413, 26857, 25881, 25349, 24736, 
    24173, 23710,
  26950, 27077, 27035, 26865, 26154, 24801, 23394, 22724, 22446, 22593, 
    22914, 23553, 24532, 25803, 26669, 27343, 26963, 26097, 25533, 24878, 
    24267, 23735,
  26829, 26977, 26980, 26818, 26151, 24854, 23478, 22765, 22470, 22584, 
    22885, 23635, 24543, 25651, 26816, 27255, 27041, 26281, 25689, 25080, 
    24278, 23747,
  26694, 26886, 26901, 26741, 26122, 24896, 23490, 22846, 22467, 22566, 
    22828, 23353, 24418, 25684, 26351, 27209, 27109, 26478, 25919, 25213, 
    24447, 23886,
  26603, 26804, 26750, 26688, 26093, 24929, 23535, 22850, 22510, 22554, 
    22825, 23559, 24412, 25696, 26491, 27182, 27311, 26617, 26040, 25391, 
    24535, 23910,
  26583, 26755, 26670, 26632, 26129, 25006, 23572, 22862, 22504, 22548, 
    22955, 23532, 24346, 25593, 26721, 27179, 27315, 26643, 26169, 25507, 
    24678, 24007,
  26626, 26750, 26719, 26657, 26142, 24993, 23592, 22925, 22530, 22607, 
    22919, 23532, 24305, 25257, 26313, 27124, 27246, 26671, 26140, 25485, 
    24664, 23971,
  26680, 26781, 26798, 26625, 26170, 25053, 23623, 22936, 22551, 22593, 
    22926, 23445, 24415, 25531, 26615, 27094, 27188, 26550, 26076, 25428, 
    24680, 24003,
  26710, 26793, 26737, 26610, 26194, 25051, 23665, 23006, 22590, 22654, 
    22881, 23491, 24391, 25342, 26416, 27046, 27226, 26685, 26276, 25577, 
    24735, 24068,
  26673, 26735, 26650, 26616, 26153, 25089, 23682, 22994, 22612, 22642, 
    22929, 23453, 24307, 25546, 26804, 27035, 27191, 26735, 26304, 25762, 
    24952, 24254,
  26561, 26596, 26579, 26560, 26125, 25080, 23693, 22987, 22623, 22661, 
    22949, 23437, 24328, 25530, 26888, 26898, 27072, 26686, 26228, 25804, 
    25010, 24315,
  26395, 26437, 26535, 26503, 26194, 25064, 23756, 23007, 22617, 22619, 
    22976, 23375, 24208, 25584, 26645, 26891, 27023, 26707, 26334, 25831, 
    25162, 24455,
  26249, 26327, 26509, 26496, 26132, 25135, 23807, 23042, 22680, 22590, 
    22974, 23416, 24256, 25479, 26401, 26878, 27050, 26735, 26360, 25851, 
    25143, 24408,
  26186, 26300, 26396, 26482, 26121, 25153, 23754, 23111, 22687, 22632, 
    22857, 23434, 24262, 25471, 26621, 26890, 27153, 26722, 26301, 25837, 
    25117, 24420,
  26211, 26344, 26388, 26485, 26158, 25186, 23812, 23098, 22699, 22646, 
    22940, 23485, 24171, 25579, 26781, 26831, 27304, 26782, 26323, 25841, 
    25186, 24419,
  26281, 26404, 26506, 26513, 26154, 25139, 23803, 23126, 22673, 22654, 
    22957, 23484, 24268, 25488, 26601, 26837, 27042, 26643, 26328, 25847, 
    25139, 24578,
  26329, 26430, 26576, 26526, 26159, 25170, 23870, 23133, 22708, 22676, 
    22896, 23338, 24396, 25399, 26944, 26920, 27114, 26675, 26204, 25715, 
    25099, 24542,
  26303, 26378, 26425, 26491, 26126, 25140, 23881, 23159, 22822, 22736, 
    22951, 23443, 24249, 25387, 26556, 26885, 27253, 26631, 26243, 25750, 
    25161, 24628,
  26193, 26253, 26391, 26427, 26147, 25186, 23877, 23178, 22742, 22678, 
    22910, 23528, 24249, 25434, 26522, 26757, 27216, 26703, 26240, 25804, 
    25166, 24708,
  26021, 26075, 26238, 26362, 26094, 25166, 23847, 23198, 22801, 22672, 
    22895, 23405, 24332, 25431, 26756, 26657, 27110, 26582, 26236, 25803, 
    25293, 24882,
  25827, 25890, 26103, 26249, 26106, 25153, 23939, 23212, 22791, 22703, 
    22978, 23443, 24265, 25515, 26299, 26476, 27101, 26587, 26234, 25839, 
    25363, 24969,
  25666, 25751, 26010, 26217, 26037, 25206, 23913, 23229, 22802, 22677, 
    22899, 23398, 24214, 25604, 26900, 26431, 26907, 26496, 26168, 25781, 
    25426, 24991,
  25619, 25729, 26037, 26192, 26060, 25139, 23900, 23217, 22802, 22735, 
    22895, 23443, 24281, 25428, 26570, 26437, 26957, 26391, 26090, 25726, 
    25363, 24971,
  25746, 25868, 26063, 26207, 26027, 25160, 23967, 23248, 22833, 22637, 
    22905, 23394, 24419, 25302, 26474, 26462, 27002, 26403, 26014, 25625, 
    25159, 24857,
  26048, 26155, 26357, 26457, 26151, 25202, 23936, 23260, 22840, 22733, 
    22919, 23418, 24309, 25532, 26453, 26644, 26984, 26359, 25916, 25564, 
    25038, 24696,
  26436, 26531, 26694, 26610, 26182, 25224, 23952, 23242, 22830, 22660, 
    22936, 23586, 24143, 25300, 26723, 26891, 26978, 26334, 25916, 25440, 
    24915, 24515,
  26790, 26899, 26744, 26646, 26249, 25296, 23981, 23271, 22801, 22727, 
    22919, 23430, 24232, 25570, 26659, 26925, 26985, 26347, 25875, 25472, 
    24871, 24541,
  27030, 27183, 26767, 26573, 26231, 25261, 23928, 23234, 22851, 22736, 
    23001, 23409, 24276, 25437, 26360, 26890, 26785, 26216, 25868, 25427, 
    24934, 24443,
  27137, 27329, 26796, 26630, 26231, 25283, 23952, 23237, 22883, 22652, 
    23037, 23419, 24141, 25424, 26844, 26879, 27021, 26344, 25888, 25464, 
    24838, 24409,
  27118, 27331, 26747, 26648, 26265, 25288, 23994, 23304, 22848, 22754, 
    22941, 23431, 24330, 25631, 26692, 26974, 27140, 26413, 25916, 25457, 
    24896, 24391,
  26976, 27176, 26779, 26719, 26234, 25302, 23966, 23267, 22927, 22745, 
    22960, 23443, 24172, 25350, 26307, 26973, 27232, 26451, 25985, 25420, 
    24992, 24453,
  26682, 26840, 26769, 26710, 26286, 25323, 23996, 23265, 22857, 22681, 
    22992, 23412, 24269, 25349, 26359, 26903, 27113, 26385, 25846, 25364, 
    24764, 24326,
  26204, 26311, 26497, 26620, 26201, 25267, 23981, 23340, 22888, 22759, 
    22939, 23457, 24223, 25260, 26600, 26766, 26835, 26225, 25713, 25214, 
    24746, 24288,
  25548, 25631, 26204, 26404, 26165, 25289, 24000, 23252, 22883, 22770, 
    22923, 23421, 24252, 25471, 26582, 26475, 26682, 25990, 25589, 25222, 
    24733, 24295,
  24792, 24877, 25756, 26046, 25996, 25232, 23985, 23321, 22919, 22725, 
    23019, 23493, 24083, 25390, 26540, 25884, 26597, 26154, 25723, 25303, 
    24727, 24282,
  24049, 24156, 25238, 25716, 25911, 25226, 23985, 23293, 22869, 22774, 
    22919, 23399, 24166, 25406, 26232, 25318, 26599, 26594, 26018, 25409, 
    24841, 24469,
  23449, 23580, 25079, 25644, 25882, 25196, 24002, 23286, 22946, 22817, 
    22963, 23431, 24273, 25328, 26585, 25064, 26679, 26846, 26325, 25578, 
    24988, 24389,
  23067, 23224, 24911, 25499, 25822, 25189, 23987, 23287, 22917, 22770, 
    23042, 23434, 24235, 25236, 26429, 24935, 26779, 26945, 26365, 25728, 
    25077, 24481,
  22937, 23097, 24792, 25451, 25797, 25176, 23971, 23290, 22895, 22757, 
    22994, 23372, 24192, 25392, 26447, 24771, 26894, 26976, 26499, 25799, 
    25031, 24512,
  23001, 23141, 24745, 25426, 25775, 25186, 23990, 23301, 22902, 22771, 
    22990, 23388, 24249, 25405, 26522, 24816, 26897, 26967, 26460, 25950, 
    25152, 24625,
  23132, 23246, 24849, 25537, 25754, 25173, 24026, 23310, 22914, 22788, 
    23048, 23385, 24149, 25489, 26434, 24966, 27021, 26994, 26459, 25874, 
    25101, 24577,
  23163, 23285, 24933, 25496, 25753, 25160, 23984, 23319, 22900, 22785, 
    22990, 23378, 24317, 25282, 26315, 25084, 26853, 26907, 26434, 25813, 
    25119, 24497,
  23019, 23168, 24860, 25433, 25718, 25135, 23972, 23266, 22951, 22799, 
    23064, 23352, 24178, 25421, 26322, 24967, 26896, 26954, 26453, 25822, 
    25087, 24431,
  22700, 22878, 24583, 25285, 25610, 25135, 23950, 23280, 22975, 22775, 
    22928, 23383, 24168, 25226, 26657, 24705, 26598, 26890, 26476, 25813, 
    25062, 24491,
  22263, 22455, 24251, 25040, 25515, 25118, 24001, 23290, 22914, 22809, 
    23029, 23507, 24313, 25317, 26571, 24427, 26313, 26826, 26424, 25865, 
    25094, 24505,
  21782, 21999, 23877, 24797, 25406, 25026, 23925, 23346, 22908, 22796, 
    22947, 23411, 24191, 25390, 26582, 24032, 26081, 26776, 26355, 25840, 
    25101, 24533,
  21328, 21590, 23699, 24662, 25315, 25037, 23983, 23342, 22938, 22862, 
    23096, 23466, 24329, 25542, 26834, 23643, 25913, 26694, 26421, 25896, 
    25088, 24485,
  20968, 21275, 23579, 24646, 25291, 24977, 23908, 23268, 22928, 22836, 
    23065, 23550, 24297, 25370, 26672, 23655, 26062, 26693, 26426, 25879, 
    25171, 24505,
  20759, 21075, 23521, 24590, 25303, 24972, 23936, 23324, 22947, 22816, 
    23006, 23517, 24181, 25412, 26692, 23589, 25997, 26741, 26488, 25891, 
    25330, 24641,
  20713, 21029, 23578, 24596, 25293, 24960, 23934, 23316, 22973, 22847, 
    23046, 23476, 24161, 25437, 26658, 23503, 25863, 26811, 26488, 26034, 
    25337, 24721,
  20811, 21117, 23812, 24691, 25315, 24931, 23904, 23269, 22992, 22886, 
    23028, 23415, 24182, 25407, 26533, 23670, 25938, 26801, 26515, 26012, 
    25326, 24842,
  21033, 21320, 23965, 24817, 25306, 24909, 23881, 23294, 22964, 22826, 
    23008, 23537, 24260, 25472, 26168, 23902, 26141, 26763, 26540, 25998, 
    25373, 24803,
  21327, 21607, 24075, 24833, 25356, 24955, 23877, 23262, 22980, 22851, 
    22982, 23518, 24371, 25521, 26656, 23998, 26119, 26738, 26513, 26012, 
    25362, 24757,
  21646, 21935, 23983, 24809, 25384, 24954, 23900, 23301, 22951, 22858, 
    23032, 23379, 24377, 25619, 26604, 23859, 25865, 26693, 26438, 26019, 
    25312, 24721,
  21961, 22241, 24125, 24875, 25343, 24877, 23854, 23268, 22975, 22868, 
    23070, 23509, 24445, 25471, 26591, 23915, 25895, 26662, 26466, 25913, 
    25332, 24709,
  22238, 22482, 24268, 24971, 25400, 24925, 23824, 23258, 22963, 22915, 
    23103, 23545, 24372, 25241, 26352, 24046, 25920, 26676, 26404, 25950, 
    25337, 24796,
  22442, 22645, 24336, 25000, 25427, 24896, 23793, 23242, 22937, 22897, 
    23086, 23508, 24276, 25376, 26560, 24111, 25925, 26703, 26449, 25944, 
    25345, 24831,
  22546, 22735, 24389, 25025, 25392, 24883, 23815, 23249, 22981, 22887, 
    23151, 23438, 24356, 25438, 26384, 24126, 25974, 26689, 26390, 25899, 
    25359, 24876,
  22521, 22729, 24293, 25027, 25385, 24831, 23809, 23260, 22983, 22845, 
    23160, 23547, 24362, 25721, 26507, 24202, 26072, 26721, 26307, 25921, 
    25270, 24799,
  22352, 22573, 24356, 25009, 25364, 24857, 23795, 23282, 22984, 22920, 
    23065, 23519, 24332, 25539, 26788, 24343, 26157, 26644, 26292, 25806, 
    25284, 24754,
  22030, 22235, 24404, 25083, 25367, 24778, 23770, 23247, 23009, 22949, 
    23077, 23594, 24334, 25592, 26737, 24460, 26300, 26610, 26310, 25859, 
    25272, 24835,
  21566, 21762, 24267, 24967, 25315, 24788, 23757, 23240, 23016, 22973, 
    23116, 23534, 24411, 25562, 26773, 24320, 26178, 26579, 26249, 25729, 
    25180, 24649,
  21061, 21287, 23897, 24851, 25309, 24768, 23772, 23277, 23003, 22937, 
    23106, 23517, 24231, 25439, 26776, 23991, 26077, 26526, 26216, 25796, 
    25129, 24626,
  20684, 20983, 23666, 24676, 25234, 24753, 23707, 23243, 22995, 22971, 
    23115, 23501, 24404, 25586, 26606, 23829, 26031, 26538, 26131, 25598, 
    25036, 24601,
  20599, 20952, 23635, 24609, 25192, 24709, 23728, 23262, 22991, 23009, 
    23137, 23486, 24543, 25632, 26583, 23719, 26004, 26457, 26123, 25584, 
    25037, 24488,
  20828, 21191, 23647, 24718, 25214, 24690, 23718, 23267, 22995, 22939, 
    23092, 23565, 24427, 25682, 26962, 23796, 25927, 26454, 26179, 25729, 
    25128, 24623,
  21269, 21589, 23954, 24867, 25257, 24687, 23689, 23214, 23016, 22976, 
    23127, 23528, 24431, 25744, 26849, 24048, 26052, 26546, 26172, 25699, 
    25090, 24585,
  21721, 22019, 24208, 24954, 25310, 24656, 23689, 23246, 23041, 22940, 
    23112, 23610, 24454, 25601, 26872, 24278, 26053, 26507, 26151, 25732, 
    25117, 24564,
  22053, 22355, 24383, 25060, 25297, 24671, 23656, 23259, 23048, 23047, 
    23077, 23626, 24548, 25794, 27125, 24475, 26153, 26504, 26149, 25716, 
    25087, 24485,
  22202, 22530, 24422, 25056, 25293, 24645, 23656, 23220, 23035, 23032, 
    23192, 23656, 24450, 25667, 26962, 24550, 26303, 26524, 26193, 25737, 
    25127, 24566,
  22232, 22546, 24321, 25067, 25242, 24552, 23661, 23227, 23043, 22981, 
    23167, 23604, 24509, 25859, 26923, 24369, 26100, 26497, 26207, 25856, 
    25097, 24668,
  22206, 22512, 24344, 25070, 25281, 24568, 23582, 23256, 23050, 23036, 
    23194, 23640, 24526, 25682, 27030, 24225, 25934, 26510, 26232, 25865, 
    25239, 24703,
  22199, 22489, 24441, 25093, 25281, 24529, 23578, 23204, 23038, 23112, 
    23264, 23719, 24619, 25890, 26960, 24267, 25991, 26500, 26234, 25823, 
    25176, 24704,
  22216, 22497, 24519, 25189, 25316, 24516, 23562, 23202, 23054, 23091, 
    23196, 23638, 24570, 25760, 27100, 24361, 26161, 26472, 26207, 25768, 
    25260, 24705,
  22246, 22513, 24596, 25169, 25224, 24514, 23546, 23228, 23050, 23031, 
    23248, 23714, 24672, 25644, 26725, 24350, 26097, 26513, 26242, 25786, 
    25184, 24640,
  22281, 22549, 24669, 25246, 25193, 24434, 23485, 23203, 23078, 23026, 
    23183, 23712, 24685, 25863, 26956, 24390, 26197, 26460, 26104, 25706, 
    25171, 24534,
  22373, 22634, 24749, 25276, 25223, 24384, 23535, 23204, 23065, 23105, 
    23201, 23695, 24636, 25766, 26918, 24603, 26360, 26446, 26048, 25657, 
    25037, 24461,
  22555, 22801, 24846, 25368, 25213, 24307, 23455, 23194, 23099, 23093, 
    23206, 23718, 24658, 26029, 26837, 24709, 26375, 26468, 26067, 25716, 
    25140, 24589,
  22837, 23057, 25065, 25400, 25210, 24317, 23466, 23223, 23080, 23045, 
    23263, 23737, 24670, 25875, 26807, 24747, 26371, 26410, 26039, 25579, 
    25033, 24496,
  23191, 23375, 25169, 25491, 25185, 24272, 23443, 23221, 23126, 23054, 
    23209, 23757, 24737, 25938, 27001, 24845, 26344, 26327, 25951, 25586, 
    24944, 24482,
  23554, 23701, 25328, 25555, 25142, 24226, 23421, 23214, 23135, 23053, 
    23282, 23832, 24915, 26225, 27140, 24850, 26307, 26296, 25960, 25481, 
    24888, 24382,
  23864, 23959, 25389, 25534, 25129, 24247, 23440, 23208, 23144, 23180, 
    23321, 23775, 24797, 26214, 27203, 24572, 26100, 26287, 25909, 25416, 
    24941, 24431,
  24088, 24121, 25332, 25511, 25054, 24217, 23401, 23197, 23114, 23147, 
    23320, 23895, 24865, 26225, 26574, 24279, 25926, 26260, 25912, 25520, 
    24893, 24520,
  24154, 24128, 25370, 25501, 25022, 24130, 23343, 23237, 23187, 23172, 
    23340, 23853, 25001, 26221, 27540, 24188, 25976, 26159, 25778, 25367, 
    24958, 24376,
  24016, 23948, 25412, 25464, 24951, 24103, 23389, 23217, 23168, 23150, 
    23348, 23964, 24876, 26200, 27019, 24104, 25784, 26071, 25724, 25289, 
    24758, 24326,
  23700, 23634, 25364, 25477, 24891, 23961, 23357, 23225, 23179, 23159, 
    23368, 23931, 25011, 26319, 27495, 24224, 25807, 26037, 25679, 25285, 
    24740, 24229,
  23544, 23469, 25446, 25477, 24843, 23975, 23293, 23232, 23160, 23137, 
    23387, 24034, 25012, 26291, 27385, 24497, 26071, 25932, 25632, 25175, 
    24601, 24029,
  27320, 27241, 27343, 26772, 25647, 24098, 22773, 22372, 22250, 22597, 
    22983, 23662, 24720, 25823, 26947, 27662, 27040, 26179, 25546, 25015, 
    24322, 23753,
  27296, 27224, 27249, 26815, 25732, 24203, 22867, 22386, 22215, 22596, 
    22970, 23749, 24837, 25713, 26815, 27688, 27304, 26248, 25665, 25078, 
    24436, 23706,
  27247, 27206, 27055, 26672, 25726, 24286, 22960, 22410, 22256, 22590, 
    22933, 23705, 24887, 25895, 26726, 27326, 27090, 26258, 25646, 25060, 
    24374, 23781,
  27185, 27189, 26945, 26623, 25750, 24393, 23012, 22514, 22334, 22639, 
    22923, 23668, 24667, 25976, 26763, 27013, 26674, 26090, 25594, 25021, 
    24406, 23612,
  27196, 27217, 26932, 26659, 25816, 24450, 23087, 22491, 22339, 22558, 
    22911, 23607, 24616, 25810, 26688, 26982, 26704, 26000, 25407, 24871, 
    24215, 23558,
  27217, 27237, 27079, 26772, 25907, 24576, 23179, 22585, 22377, 22587, 
    22901, 23629, 24516, 25823, 26666, 27204, 26921, 25924, 25361, 24755, 
    24145, 23517,
  27622, 27572, 27244, 26785, 25898, 24557, 23183, 22479, 22343, 22542, 
    22939, 23543, 24490, 25614, 26982, 27481, 26479, 25418, 25021, 24556, 
    24086, 23477,
  27593, 27563, 27254, 26856, 25975, 24667, 23227, 22547, 22355, 22550, 
    22942, 23589, 24541, 25818, 26571, 27557, 26423, 25468, 25000, 24556, 
    24149, 23564,
  27144, 27221, 27126, 26932, 26115, 24760, 23334, 22700, 22448, 22614, 
    22956, 23596, 24576, 25622, 26985, 27417, 26770, 25813, 25258, 24816, 
    24261, 23584,
  27088, 27177, 27060, 26939, 26190, 24776, 23399, 22688, 22436, 22579, 
    22967, 23541, 24630, 25642, 26540, 27453, 27021, 26176, 25524, 25009, 
    24248, 23786,
  26997, 27084, 27079, 26908, 26159, 24821, 23376, 22776, 22451, 22501, 
    22896, 23564, 24485, 25731, 26522, 27413, 27107, 26328, 25679, 25157, 
    24354, 23737,
  26867, 26985, 27026, 26898, 26194, 24879, 23457, 22812, 22508, 22564, 
    22860, 23521, 24449, 25640, 26461, 27354, 27160, 26462, 25871, 25229, 
    24468, 23924,
  26714, 26897, 26878, 26763, 26124, 24919, 23521, 22821, 22502, 22544, 
    22920, 23470, 24351, 25570, 26608, 27338, 27252, 26500, 26006, 25399, 
    24580, 23962,
  26599, 26805, 26782, 26700, 26096, 24961, 23510, 22852, 22486, 22649, 
    22903, 23460, 24433, 25769, 26703, 27244, 27330, 26726, 26119, 25534, 
    24731, 24013,
  26551, 26733, 26703, 26676, 26134, 24999, 23582, 22855, 22532, 22611, 
    22885, 23501, 24437, 25621, 26910, 27178, 27272, 26703, 26150, 25512, 
    24746, 24042,
  26571, 26706, 26748, 26663, 26145, 25000, 23622, 22904, 22550, 22525, 
    22969, 23439, 24342, 25679, 26508, 27123, 27271, 26635, 26142, 25559, 
    24688, 23913,
  26623, 26729, 26743, 26667, 26092, 24993, 23619, 22917, 22539, 22625, 
    22848, 23407, 24417, 25518, 26361, 27106, 27189, 26694, 26190, 25682, 
    24762, 24099,
  26679, 26757, 26707, 26628, 26119, 25024, 23700, 22982, 22629, 22637, 
    22950, 23403, 24504, 25491, 26572, 27092, 27196, 26744, 26328, 25750, 
    24939, 24278,
  26689, 26740, 26659, 26563, 26146, 25076, 23716, 23014, 22629, 22542, 
    22885, 23441, 24277, 25546, 26809, 27005, 27179, 26743, 26369, 25824, 
    25122, 24370,
  26635, 26664, 26631, 26560, 26182, 25076, 23747, 22996, 22617, 22670, 
    22887, 23425, 24453, 25214, 26535, 26947, 26991, 26686, 26313, 25854, 
    25117, 24338,
  26527, 26580, 26627, 26570, 26168, 25132, 23726, 23056, 22660, 22649, 
    22854, 23426, 24401, 25552, 26576, 26947, 27099, 26715, 26287, 25887, 
    25174, 24351,
  26432, 26540, 26547, 26566, 26120, 25123, 23789, 23070, 22679, 22607, 
    22941, 23426, 24364, 25565, 26809, 26929, 27051, 26713, 26281, 25813, 
    25174, 24297,
  26405, 26558, 26458, 26543, 26129, 25104, 23754, 23054, 22693, 22673, 
    22850, 23472, 24210, 25467, 26773, 26933, 27160, 26759, 26255, 25849, 
    25243, 24376,
  26448, 26615, 26491, 26505, 26129, 25131, 23836, 23127, 22626, 22634, 
    22864, 23458, 24271, 25596, 26372, 26904, 27068, 26710, 26319, 25866, 
    25249, 24468,
  26523, 26665, 26608, 26584, 26123, 25129, 23798, 23122, 22710, 22619, 
    22851, 23406, 24324, 25511, 26670, 26961, 26986, 26600, 26151, 25822, 
    25215, 24647,
  26569, 26680, 26572, 26547, 26147, 25149, 23838, 23176, 22736, 22621, 
    22912, 23455, 24304, 25476, 26824, 26972, 27114, 26619, 26200, 25752, 
    25257, 24631,
  26536, 26629, 26471, 26531, 26128, 25155, 23859, 23163, 22724, 22607, 
    22882, 23372, 24224, 25599, 26337, 26841, 27122, 26597, 26182, 25850, 
    25337, 24811,
  26409, 26505, 26385, 26434, 26154, 25154, 23900, 23159, 22733, 22667, 
    22849, 23467, 24418, 25427, 26574, 26654, 26836, 26552, 26249, 25829, 
    25331, 24811,
  26201, 26300, 26387, 26415, 26090, 25190, 23898, 23178, 22800, 22620, 
    22919, 23408, 24187, 25184, 26711, 26639, 26706, 26424, 26114, 25746, 
    25394, 24945,
  25937, 26040, 26459, 26377, 26109, 25185, 23921, 23175, 22843, 22683, 
    22905, 23432, 24311, 25255, 26279, 26653, 26866, 26428, 26091, 25857, 
    25349, 24918,
  25667, 25779, 26318, 26364, 26137, 25160, 23957, 23202, 22810, 22680, 
    22928, 23374, 24157, 25357, 26381, 26603, 26939, 26503, 26081, 25756, 
    25425, 25006,
  25485, 25609, 26000, 26185, 26039, 25137, 23937, 23251, 22801, 22680, 
    22838, 23442, 24135, 25249, 26839, 26413, 26932, 26494, 26045, 25694, 
    25330, 24946,
  25486, 25607, 25856, 26099, 26044, 25181, 23901, 23208, 22838, 22660, 
    22846, 23357, 24130, 25185, 26835, 26254, 26859, 26338, 25913, 25494, 
    25113, 24711,
  25710, 25803, 26113, 26267, 26100, 25218, 23931, 23276, 22843, 22676, 
    22872, 23479, 24318, 25292, 26663, 26436, 26816, 26279, 25829, 25439, 
    24979, 24497,
  26098, 26168, 26551, 26515, 26171, 25287, 23986, 23246, 22832, 22698, 
    22866, 23431, 24199, 25309, 26252, 26813, 26717, 26116, 25725, 25458, 
    24927, 24458,
  26527, 26600, 26737, 26634, 26231, 25243, 23977, 23273, 22834, 22799, 
    22952, 23484, 24175, 25526, 26616, 26932, 26744, 26203, 25794, 25347, 
    24895, 24456,
  26880, 26983, 26735, 26658, 26222, 25262, 23969, 23224, 22818, 22701, 
    22901, 23359, 24181, 25428, 26099, 26894, 26835, 26209, 25774, 25333, 
    24742, 24338,
  27080, 27209, 26788, 26680, 26224, 25245, 23947, 23276, 22853, 22716, 
    22929, 23356, 24225, 25363, 26572, 26933, 26990, 26294, 25774, 25302, 
    24812, 24365,
  27081, 27235, 26803, 26688, 26221, 25295, 24004, 23324, 22847, 22686, 
    22885, 23464, 24226, 25179, 26218, 26970, 26822, 26175, 25676, 25264, 
    24786, 24420,
  26869, 27029, 26783, 26686, 26265, 25284, 24010, 23277, 22876, 22690, 
    22742, 23358, 24151, 25492, 26559, 26930, 26654, 26032, 25607, 25189, 
    24800, 24241,
  26426, 26571, 26688, 26576, 26270, 25311, 24033, 23299, 22912, 22707, 
    22893, 23425, 24228, 25039, 26591, 26876, 26591, 25972, 25558, 25158, 
    24635, 24214,
  25752, 25866, 26318, 26392, 26128, 25251, 23993, 23311, 22846, 22728, 
    23003, 23458, 24200, 25180, 26404, 26573, 26644, 26088, 25666, 25245, 
    24763, 24303,
  24891, 24996, 25812, 26098, 26024, 25239, 24013, 23327, 22850, 22756, 
    22958, 23363, 24318, 25264, 26582, 26035, 26814, 26438, 25875, 25408, 
    24808, 24298,
  23974, 24089, 25237, 25747, 25875, 25270, 23978, 23296, 22886, 22716, 
    22874, 23415, 24270, 25413, 26459, 25332, 26672, 26595, 26133, 25589, 
    24981, 24385,
  23162, 23303, 24858, 25535, 25811, 25188, 23967, 23312, 22865, 22676, 
    22858, 23354, 24348, 25492, 26461, 24851, 26629, 26869, 26276, 25700, 
    25031, 24438,
  22610, 22776, 24751, 25462, 25778, 25220, 24012, 23347, 22934, 22748, 
    22942, 23416, 24149, 25306, 26880, 24745, 26874, 26910, 26376, 25788, 
    25127, 24504,
  22369, 22559, 24572, 25353, 25747, 25154, 24020, 23369, 22910, 22707, 
    22881, 23475, 24250, 25225, 26717, 24560, 26754, 26938, 26403, 25834, 
    25140, 24556,
  22416, 22599, 24466, 25253, 25633, 25151, 23976, 23371, 22914, 22751, 
    22881, 23396, 24332, 25427, 26196, 24241, 26408, 26890, 26397, 25799, 
    25144, 24454,
  22621, 22768, 24441, 25210, 25581, 25084, 23951, 23296, 22905, 22754, 
    22937, 23505, 24259, 25305, 26514, 24124, 26050, 26794, 26325, 25788, 
    25100, 24507,
  22802, 22906, 24548, 25215, 25604, 25071, 23982, 23327, 22896, 22825, 
    22912, 23442, 24284, 25070, 26526, 24137, 25954, 26754, 26344, 25849, 
    25010, 24492,
  22775, 22878, 24472, 25182, 25566, 25075, 23973, 23320, 22916, 22776, 
    22944, 23427, 24317, 25437, 26649, 24175, 25962, 26713, 26326, 25738, 
    24927, 24466,
  22494, 22625, 24310, 25071, 25497, 25075, 23964, 23314, 22876, 22799, 
    23042, 23393, 24246, 25533, 26669, 24027, 25899, 26666, 26351, 25822, 
    25060, 24393,
  22026, 22188, 24046, 24882, 25399, 25011, 23977, 23291, 22924, 22781, 
    23004, 23503, 24308, 25464, 26553, 23738, 25763, 26667, 26326, 25837, 
    25163, 24454,
  21488, 21664, 23739, 24684, 25371, 25001, 23923, 23304, 22934, 22795, 
    22976, 23447, 24256, 25229, 26507, 23468, 25709, 26669, 26419, 25778, 
    25125, 24526,
  20990, 21188, 23446, 24486, 25205, 25008, 23958, 23274, 22899, 22791, 
    23087, 23360, 24346, 25276, 26413, 23164, 25721, 26669, 26398, 25871, 
    25189, 24595,
  20606, 20844, 23329, 24460, 25163, 24951, 23933, 23329, 22972, 22818, 
    22974, 23416, 24323, 25463, 26848, 23096, 25732, 26766, 26457, 26020, 
    25285, 24615,
  20390, 20670, 23415, 24446, 25225, 24930, 23962, 23293, 22989, 22836, 
    23040, 23436, 24392, 25516, 26438, 23266, 25913, 26772, 26428, 26060, 
    25335, 24722,
  20378, 20668, 23375, 24473, 25239, 24973, 23949, 23308, 22946, 22782, 
    22939, 23459, 24262, 25321, 26558, 23301, 25910, 26763, 26429, 25966, 
    25336, 24716,
  20549, 20841, 23574, 24562, 25278, 24939, 23930, 23321, 22984, 22847, 
    22926, 23499, 24299, 25307, 26378, 23496, 25951, 26775, 26442, 26109, 
    25350, 24797,
  20840, 21128, 23876, 24766, 25342, 24924, 23886, 23339, 22918, 22828, 
    23126, 23507, 24386, 25357, 26551, 23847, 26182, 26808, 26516, 26092, 
    25402, 24831,
  21196, 21470, 24035, 24811, 25328, 24938, 23905, 23316, 22968, 22814, 
    23075, 23351, 24282, 25342, 26806, 24029, 26122, 26763, 26494, 26040, 
    25442, 24899,
  21556, 21815, 24053, 24802, 25333, 24926, 23884, 23278, 22983, 22874, 
    23007, 23390, 24193, 25349, 26369, 23941, 25889, 26673, 26440, 26035, 
    25392, 24940,
  21879, 22130, 24102, 24861, 25349, 24912, 23867, 23256, 22939, 22852, 
    23056, 23434, 24354, 25638, 26460, 23902, 25859, 26686, 26385, 26094, 
    25406, 24817,
  22159, 22384, 24212, 24972, 25331, 24895, 23864, 23240, 22883, 22863, 
    22999, 23505, 24336, 25431, 26660, 23955, 25958, 26704, 26461, 26025, 
    25368, 24918,
  22385, 22573, 24279, 25010, 25353, 24890, 23844, 23272, 22963, 22924, 
    23135, 23515, 24416, 25523, 26466, 23919, 25802, 26669, 26351, 25974, 
    25387, 24920,
  22546, 22695, 24223, 25004, 25380, 24887, 23851, 23279, 22984, 22895, 
    23136, 23483, 24268, 25709, 26649, 23882, 25770, 26669, 26375, 25912, 
    25387, 24812,
  22610, 22746, 24288, 25024, 25371, 24912, 23836, 23257, 22992, 22911, 
    23055, 23512, 24334, 25391, 26633, 23962, 25856, 26639, 26385, 25893, 
    25282, 24832,
  22529, 22688, 24276, 25056, 25399, 24833, 23807, 23297, 22935, 22817, 
    23129, 23639, 24342, 25505, 26869, 24131, 25949, 26620, 26240, 25802, 
    25231, 24795,
  22278, 22471, 24329, 25044, 25353, 24850, 23832, 23271, 22998, 22893, 
    23118, 23606, 24416, 25422, 26522, 24334, 26057, 26578, 26219, 25781, 
    25168, 24668,
  21870, 22078, 24399, 25084, 25369, 24827, 23797, 23252, 23006, 22923, 
    23052, 23533, 24418, 25682, 26918, 24506, 26263, 26466, 26147, 25665, 
    25112, 24596,
  21356, 21580, 24161, 24958, 25318, 24815, 23732, 23244, 22978, 22921, 
    23152, 23524, 24361, 25835, 26876, 24414, 26235, 26507, 26162, 25637, 
    25070, 24564,
  20868, 21138, 23682, 24683, 25245, 24730, 23771, 23229, 23020, 22950, 
    23104, 23475, 24357, 25775, 26690, 23897, 26027, 26520, 26094, 25709, 
    25026, 24501,
  20576, 20924, 23413, 24556, 25202, 24690, 23769, 23224, 22968, 22910, 
    23176, 23502, 24401, 25521, 26646, 23725, 26025, 26424, 26086, 25622, 
    25073, 24617,
  20609, 21001, 23570, 24642, 25172, 24727, 23745, 23228, 23016, 22929, 
    23115, 23601, 24306, 25570, 26572, 23787, 26010, 26529, 26167, 25738, 
    25125, 24544,
  20941, 21317, 23774, 24768, 25216, 24677, 23665, 23242, 22970, 22953, 
    23110, 23586, 24384, 25516, 26580, 23951, 25971, 26569, 26201, 25716, 
    25171, 24659,
  21438, 21743, 24105, 24931, 25278, 24675, 23699, 23262, 23016, 22942, 
    23089, 23521, 24468, 25769, 26611, 24178, 26096, 26532, 26154, 25735, 
    25217, 24621,
  21907, 22177, 24382, 25074, 25306, 24671, 23667, 23248, 22976, 23004, 
    23105, 23697, 24505, 25535, 26457, 24468, 26109, 26479, 26113, 25688, 
    25180, 24586,
  22237, 22513, 24533, 25161, 25340, 24637, 23680, 23243, 23040, 22959, 
    23163, 23692, 24469, 25682, 26976, 24649, 26259, 26476, 26110, 25722, 
    25054, 24594,
  22376, 22690, 24476, 25168, 25320, 24632, 23669, 23225, 23061, 23009, 
    23195, 23600, 24602, 25809, 27060, 24593, 26259, 26517, 26174, 25710, 
    25190, 24528,
  22391, 22698, 24411, 25125, 25273, 24624, 23670, 23282, 23048, 23005, 
    23188, 23729, 24567, 25729, 26588, 24289, 25982, 26504, 26176, 25732, 
    25216, 24570,
  22345, 22640, 24329, 25053, 25246, 24583, 23617, 23237, 23082, 22959, 
    23235, 23666, 24499, 25545, 26784, 24212, 25953, 26497, 26199, 25838, 
    25251, 24737,
  22316, 22585, 24482, 25114, 25189, 24522, 23584, 23227, 23066, 23043, 
    23151, 23707, 24596, 25751, 26828, 24374, 26135, 26485, 26195, 25804, 
    25271, 24726,
  22305, 22567, 24588, 25171, 25272, 24515, 23579, 23216, 23056, 23045, 
    23109, 23641, 24503, 25838, 26807, 24529, 26212, 26479, 26155, 25731, 
    25207, 24647,
  22301, 22566, 24647, 25276, 25252, 24481, 23587, 23203, 23131, 23031, 
    23214, 23679, 24531, 26053, 26806, 24546, 26222, 26463, 26120, 25600, 
    25093, 24575,
  22294, 22589, 24733, 25287, 25198, 24425, 23530, 23196, 23077, 23029, 
    23204, 23758, 24539, 25988, 27053, 24570, 26222, 26424, 26079, 25704, 
    25062, 24603,
  22347, 22659, 24819, 25301, 25220, 24413, 23531, 23215, 23141, 23083, 
    23245, 23685, 24689, 26047, 27045, 24651, 26354, 26468, 26078, 25693, 
    25029, 24511,
  22502, 22810, 24918, 25348, 25238, 24415, 23482, 23275, 23107, 23069, 
    23266, 23749, 24689, 25772, 26984, 24746, 26381, 26425, 26097, 25654, 
    25151, 24571,
  22777, 23055, 25056, 25417, 25155, 24327, 23462, 23222, 23064, 23087, 
    23247, 23860, 24596, 25917, 27010, 24782, 26409, 26360, 25985, 25604, 
    24993, 24371,
  23142, 23370, 25183, 25482, 25159, 24305, 23498, 23258, 23099, 23090, 
    23304, 23737, 24781, 25911, 27006, 24900, 26432, 26320, 25940, 25504, 
    24911, 24411,
  23527, 23703, 25344, 25514, 25147, 24265, 23434, 23210, 23137, 23105, 
    23348, 23765, 24732, 26159, 27187, 24904, 26365, 26288, 25893, 25499, 
    24855, 24311,
  23857, 23971, 25382, 25533, 25138, 24234, 23450, 23222, 23155, 23120, 
    23308, 23834, 24697, 26135, 27103, 24674, 26057, 26237, 25884, 25434, 
    24908, 24446,
  24090, 24140, 25389, 25550, 25020, 24166, 23421, 23211, 23171, 23110, 
    23246, 23900, 24854, 25910, 26907, 24299, 25890, 26289, 25928, 25514, 
    25018, 24569,
  24157, 24150, 25336, 25505, 25033, 24131, 23380, 23230, 23167, 23140, 
    23343, 23874, 24776, 26118, 27457, 24030, 25846, 26267, 25891, 25516, 
    24950, 24552,
  24024, 23975, 25344, 25447, 24930, 24071, 23395, 23243, 23167, 23141, 
    23472, 23950, 24914, 26244, 27241, 23793, 25647, 26150, 25762, 25320, 
    24909, 24395,
  23720, 23667, 25385, 25411, 24896, 23991, 23356, 23217, 23182, 23182, 
    23423, 23942, 24912, 26132, 27319, 23902, 25670, 26015, 25648, 25242, 
    24752, 24318,
  23570, 23505, 25404, 25390, 24834, 23926, 23334, 23248, 23162, 23143, 
    23368, 24022, 24947, 26400, 27282, 24199, 25922, 25875, 25545, 25125, 
    24606, 24085 ;

 CLW =
  0, 0, 0, 0, 0, 0, 0, 0, 1, 25, 0, 0, 0, 0, 49, 36, 39, 20, 2, 3, 23, 30, 
    30, 39, 40, 34, 31, 29, 33, 39, 44, 40, 45, 61, 59, 52, 41, 32, 40, 36, 
    34, 19, 7, 10, 13, 8, 1, 8, 15, 0, 1, 4, 4, 4, 5, 5, 5, 7, 5, 0, 0, 0, 4, 
    3, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 2, 1, 2, 6, 5, 2, 0, 
    0, 1, 5, 5, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 2, 14, 0, 0, 0, 0, 0, 53, 51, 31, 31, 27, 34, 33, 47, 
    52, 57, 38, 40, 33, 39, 33, 38, 37, 38, 36, 37, 34, 50, 49, 59, 47, 36, 
    27, 23, 8, 6, 6, 7, 10, 7, 3, 1, 2, 2, 3, 3, 5, 3, 3, 5, 11, 9, 0, 0, 0, 
    2, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 2, 2, 1, 2, 5, 6, 4, 0, 
    0, 2, 5, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 1, 23, 0, 0, 0, 0, 0, 54, 36, 66, 41, 32, 37, 28, 32, 33, 
    33, 32, 41, 51, 39, 38, 31, 9, 11, 17, 29, 36, 35, 34, 43, 36, 43, 39, 
    26, 24, 19, 9, 7, 6, 9, 10, 5, 1, 3, 3, 3, 4, 6, 3, 1, 3, 13, 13, 6, 0, 
    0, 2, 1, 1, 3, 2, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 0, 1, 5, 6, 1, 
    1, 0, 0, 1, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 1, 13, 36, 0, 0, 0, 0, 39, 37, 34, 38, 40, 44, 42, 33, 32, 
    44, 37, 44, 44, 38, 30, 48, 12, 25, 30, 36, 24, 39, 42, 39, 28, 28, 31, 
    33, 29, 26, 10, 7, 6, 9, 15, 21, 11, 5, 3, 2, 8, 5, 4, 4, 2, 2, 9, 12, 8, 
    0, 0, 1, 1, 1, 3, 0, 0, 0, 0, 0, 0, 1, 1, 2, 2, 2, 0, 0, 0, 0, 0, 2, 6, 
    2, 1, 1, 1, 2, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 5, 17, 22, 0, 0, 0, 0, 54, 24, 26, 44, 41, 40, 34, 34, 37, 
    58, 109, 56, 37, 53, 45, 39, 12, 10, 8, 7, 12, 33, 16, 26, 14, 11, 24, 
    26, 25, 6, 3, 3, 4, 14, 32, 10, 8, 9, 15, 13, 5, 5, 5, 2, 5, 4, 5, 9, 9, 
    0, 0, 1, 1, 2, 2, 0, 0, 0, 0, 1, 1, 1, 1, 2, 4, 1, 0, 0, 0, 0, 0, 0, 3, 
    2, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0,
  0, 3, 5, 1, 12, 1, 13, 0, 0, 0, 41, 107, 61, 41, 31, 32, 38, 33, 28, 31, 
    34, 59, 89, 35, 25, 36, 35, 40, 10, 7, 8, 6, 11, 13, 14, 28, 28, 10, 21, 
    26, 25, 6, 3, 4, 17, 7, 8, 6, 22, 33, 32, 8, 6, 3, 2, 6, 7, 7, 6, 11, 0, 
    0, 0, 1, 1, 1, 0, 0, 0, 0, 0, 2, 1, 0, 1, 3, 5, 2, 1, 0, 0, 0, 0, 0, 2, 
    3, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0,
  9, 19, 17, 17, 19, 11, 44, 0, 0, 38, 29, 67, 57, 30, 28, 35, 42, 30, 30, 
    66, 86, 71, 32, 45, 38, 31, 15, 24, 5, 4, 7, 8, 31, 38, 39, 33, 23, 11, 
    29, 28, 26, 15, 45, 71, 56, 55, 41, 23, 11, 8, 9, 5, 3, 1, 6, 4, 7, 10, 
    15, 8, 0, 0, 0, 1, 2, 1, 0, 0, 0, 0, 2, 1, 0, 0, 0, 3, 5, 4, 1, 1, 2, 0, 
    0, 2, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  7, 15, 23, 23, 13, 51, 0, 0, 0, 32, 40, 37, 28, 4, 20, 25, 6, 25, 32, 65, 
    55, 41, 33, 35, 33, 8, 33, 29, 6, 7, 9, 8, 20, 38, 36, 32, 35, 24, 22, 
    28, 26, 77, 88, 82, 66, 53, 53, 29, 5, 5, 7, 3, 3, 2, 5, 7, 12, 17, 11, 
    1, 0, 0, 1, 2, 1, 1, 0, 0, 0, 1, 1, 0, 0, 0, 1, 2, 5, 4, 3, 1, 2, 2, 1, 
    1, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0,
  14, 5, 15, 22, 33, 0, 0, 65, 28, 10, 19, 24, 30, 6, 3, 8, 37, 32, 40, 100, 
    45, 37, 30, 33, 39, 12, 87, 31, 4, 5, 8, 6, 20, 34, 43, 39, 93, 76, 32, 
    66, 90, 69, 29, 30, 30, 29, 12, 6, 4, 2, 4, 3, 7, 6, 6, 10, 14, 5, 0, 0, 
    1, 3, 2, 1, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 1, 1, 2, 2, 3, 2, 2, 2, 1, 1, 
    1, 1, 1, 2, 4, 0, 0, 0, 0, 0, 0, 0,
  8, 3, 17, 31, 76, 0, 36, 9, 2, 3, 15, 29, 27, 4, 6, 11, 30, 11, 23, 30, 29, 
    13, 35, 32, 9, 26, 31, 4, 4, 5, 5, 11, 14, 11, 11, 21, 60, 31, 18, 32, 
    43, 7, 43, 34, 14, 9, 6, 3, 5, 5, 4, 8, 11, 10, 1, 11, 13, 2, 0, 0, 1, 3, 
    2, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 2, 2, 1, 1, 0, 1, 1, 1, 1, 1, 
    1, 2, 0, 0, 0, 0, 0, 0, 0, 0,
  7, 6, 17, 49, 86, 28, 5, 1, 21, 24, 26, 28, 31, 6, 7, 14, 29, 14, 30, 34, 
    32, 41, 26, 6, 37, 28, 7, 6, 8, 6, 13, 11, 7, 9, 13, 24, 32, 9, 6, 5, 7, 
    35, 26, 20, 6, 3, 1, 0, 0, 1, 5, 2, 1, 0, 3, 0, 1, 0, 0, 1, 2, 2, 1, 0, 
    0, 0, 0, 0, 0, 2, 2, 2, 1, 1, 1, 1, 1, 1, 1, 1, 0, 1, 1, 1, 1, 2, 2, 2, 
    4, 0, 0, 0, 0, 0, 0, 0,
  14, 3, 9, 35, 30, 10, 0, 0, 26, 27, 25, 28, 9, 6, 8, 25, 35, 19, 15, 35, 
    28, 40, 25, 36, 45, 11, 7, 30, 36, 31, 19, 12, 8, 24, 39, 42, 28, 7, 34, 
    41, 46, 37, 13, 8, 3, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 2, 1, 
    0, 0, 0, 0, 0, 0, 0, 4, 4, 1, 1, 1, 1, 1, 2, 2, 1, 0, 0, 1, 1, 1, 2, 2, 
    2, 3, 3, 0, 0, 0, 0, 0, 0, 0 ;

 ChanSel =
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1 ;

 ChiSqr =
  0.1008461, 0.1342951, 0.2309889, 0.09135432, 0.08736515, 0.08311268, 
    0.118963, 0.499799, 0.4415751, 0.4981582, 0.1511773, 0.7385971, 0.711108, 
    0.600167, 0.4987307, 0.8511323, 0.6766284, 0.4243806, 0.5470757, 
    0.6629881, 0.1565461, 0.187768, 0.1674572, 0.954457, 0.1291059, 
    0.2078876, 0.1201, 0.1122698, 0.1116915, 0.2485472, 0.2671911, 0.2770049, 
    0.828739, 0.4475992, 0.199902, 0.4642757, 0.4300698, 0.7745846, 0.264123, 
    0.1750679, 0.1065845, 0.8190032, 0.6477903, 0.4421234, 0.6562275, 
    0.8462268, 1.84764, 1.084516, 0.5194832, 0.1216637, 2.061218, 0.3077135, 
    0.5300809, 0.3197876, 0.9410091, 0.3619125, 0.4276822, 0.8581687, 
    0.6692483, 0.6590104, 1.379585, 0.9880861, 0.619318, 0.506291, 0.6069245, 
    0.5390903, 0.4176021, 0.3178004, 0.5825225, 0.789907, 0.5974104, 
    0.6745406, 0.3992053, 0.923258, 0.8661819, 0.6943033, 0.8706642, 
    0.7264254, 0.5447694, 0.4560589, 0.5488386, 0.7926893, 0.4617552, 
    0.1288275, 0.07362142, 0.3113467, 0.8061541, 0.8756009, 0.817432, 
    0.6832917, 0.659427, 0.1741704, 0.1332782, 0.1986117, 0.2875583, 0.6638222,
  0.1236612, 0.1425509, 0.2550566, 0.07536855, 0.1188622, 0.08682251, 
    0.6298522, 0.5764285, 0.6855903, 0.4251214, 0.6525679, 0.3608646, 
    0.6535135, 0.9649411, 0.4353254, 0.8883732, 1.224629, 0.536883, 
    0.1185779, 0.8719167, 0.1934141, 0.8087686, 0.8578683, 0.9650786, 
    0.4514389, 0.2127961, 0.1073586, 0.1010381, 0.4867712, 0.8265147, 
    0.1405066, 0.2986663, 0.5613249, 0.4642355, 0.3205554, 0.5799623, 
    0.5322936, 0.9683701, 0.6033162, 0.2013655, 0.4421514, 0.5185236, 
    0.3749774, 0.4385787, 0.4794968, 0.4483963, 0.9897857, 0.5733235, 
    0.6496623, 0.2993832, 0.7367212, 0.6291794, 0.3191618, 0.1929728, 
    0.2950524, 0.7753845, 0.4740658, 0.4261971, 0.6600646, 0.7963629, 
    0.8127527, 1.372007, 0.9073994, 0.755116, 0.7040939, 0.409826, 0.3393357, 
    0.533318, 0.6025077, 0.9014, 0.9402861, 0.9991844, 0.8641174, 0.6788228, 
    0.6279678, 0.5397745, 0.6688898, 0.5958757, 0.672718, 0.8621103, 
    0.6551194, 0.7613919, 0.3399222, 0.05636168, 0.09935586, 0.3048741, 
    0.7953712, 0.4459568, 0.59142, 0.4065113, 0.2517513, 0.3235914, 
    0.2231312, 0.149572, 0.2901628, 0.262194,
  0.09335696, 0.1062689, 0.1200924, 0.0835233, 0.6037627, 0.6757448, 
    0.2109554, 0.3692551, 0.4004562, 0.739179, 0.6502189, 0.7833443, 
    0.5611867, 0.2995979, 1.358496, 0.93599, 0.880371, 0.3520434, 0.3668915, 
    0.1613831, 0.1363588, 0.119173, 0.17203, 0.2978281, 0.5591577, 0.3360626, 
    0.1079886, 0.1148169, 0.4657358, 0.7766832, 0.4979548, 0.6759121, 
    0.9366003, 0.2909121, 0.154625, 0.1367855, 0.2566204, 0.488337, 
    0.2398358, 0.5305606, 0.2187453, 0.8613635, 0.5328675, 0.4155954, 
    0.8443223, 0.8620353, 0.7848024, 0.8582613, 0.3313267, 0.3093867, 
    0.652791, 0.3497347, 0.5365789, 0.6232036, 0.5299205, 0.554284, 
    0.4248798, 0.3046891, 0.6445318, 0.5667638, 1.386946, 1.336446, 
    0.9883173, 0.8145404, 0.6751265, 0.4710908, 0.3101453, 0.2585951, 
    0.7304912, 0.4674543, 0.7656512, 0.615268, 0.7623305, 0.4779314, 
    0.592528, 0.3899044, 0.5694283, 0.8576469, 0.9024996, 0.891897, 
    0.9079936, 0.8325374, 0.2860918, 0.1484248, 0.3241497, 0.4399716, 
    0.7209734, 0.2827065, 0.1059716, 0.6534167, 0.1876756, 0.1455703, 
    0.1532021, 0.09721129, 0.2432538, 0.2086882,
  0.07075233, 0.9274029, 0.7985702, 0.8639729, 0.1453608, 0.2938125, 
    0.300325, 0.3319083, 0.2637465, 0.4417728, 0.7856153, 0.2392074, 
    0.4558704, 0.457949, 0.5115976, 0.8235006, 0.9406362, 0.7517352, 
    0.5400072, 0.2476903, 0.2737382, 0.4654588, 0.4651422, 0.8215367, 
    0.4576702, 0.5224178, 0.8369255, 0.1352868, 0.7012119, 0.3236287, 
    0.6046183, 0.8120943, 0.554196, 0.1271312, 0.2264372, 0.3536027, 
    0.5452742, 0.3051419, 0.2637131, 0.5907456, 0.511728, 0.9562442, 
    0.2949426, 0.337179, 0.3209908, 0.2802465, 0.3505244, 0.4625541, 
    0.3767924, 0.3016784, 0.3697577, 0.1316959, 0.3845473, 0.5486327, 
    0.5306692, 0.7328739, 0.8578034, 0.410797, 0.4961954, 0.9123142, 
    0.9970488, 0.8984271, 0.9844059, 0.8912315, 0.6229029, 0.4189267, 
    0.2180947, 0.7124293, 0.9206261, 0.4784121, 0.8041344, 0.8228258, 
    0.6270036, 0.304121, 0.3824639, 0.3004784, 0.3486047, 0.5332738, 
    0.8124743, 0.8090023, 0.6948856, 0.5825896, 0.07218481, 0.1523851, 
    0.23725, 0.3558671, 0.83801, 0.5264258, 0.7016711, 0.4598041, 0.3099987, 
    0.1221491, 0.3094735, 0.2253319, 0.2798543, 0.2084711,
  0.2258907, 0.1362204, 0.1052978, 0.4004489, 0.2595983, 0.5350647, 
    0.5975784, 0.925581, 0.8148518, 0.9908801, 0.4931153, 0.2913288, 
    0.3442559, 0.2486092, 0.1565728, 0.8986811, 1.731605, 0.9730593, 
    0.2468665, 0.7974541, 0.1870804, 0.7453068, 0.8619364, 0.2988765, 
    0.187758, 0.842362, 0.1877807, 0.2262029, 0.9841524, 0.9583538, 
    0.1437517, 0.2905164, 0.4492402, 0.2278522, 0.5743654, 0.3403841, 
    0.6965695, 0.9676022, 0.3099746, 0.19829, 0.3969177, 0.8749074, 
    0.4596163, 0.7498124, 0.3936078, 0.25582, 0.6925448, 0.1826489, 
    0.2001127, 0.2406278, 0.3580397, 0.4376269, 0.6333528, 0.3539843, 
    0.6890325, 0.7550589, 0.3809596, 0.2852807, 0.3006609, 0.4119602, 
    0.9398786, 0.8991441, 1.286627, 0.657189, 0.6784174, 0.2191618, 
    0.3392338, 0.66907, 0.346205, 0.7239518, 0.6312996, 0.2968616, 0.2767024, 
    0.489678, 0.4291223, 0.2517892, 0.3267455, 0.687529, 0.766411, 0.9685459, 
    0.7613796, 0.2496623, 0.2085657, 0.1021168, 0.2732655, 0.351776, 
    0.6519814, 0.5683877, 0.6563033, 0.2656189, 0.2562587, 0.2311982, 
    0.2098379, 0.1381075, 0.117891, 0.187325,
  0.6138157, 0.6074043, 0.8834629, 0.6020501, 0.140472, 0.9009735, 0.499988, 
    0.2529559, 0.6483934, 0.2662542, 0.2537729, 1.069554, 0.321454, 
    0.5637789, 0.6038248, 4.830637, 0.6492585, 0.2568048, 0.1731966, 
    0.08867583, 0.1033527, 0.5075077, 0.5012941, 0.5299752, 0.645685, 
    0.7369583, 0.193428, 0.6328286, 0.6351323, 0.3123596, 0.3400117, 
    0.1769601, 0.4742481, 0.5664756, 0.7555686, 0.3833653, 0.6387357, 
    0.9422989, 0.4368945, 0.2572627, 0.3508787, 0.7257026, 0.9345154, 
    0.2894699, 0.231186, 0.5391884, 0.7742103, 0.811534, 0.4676085, 
    0.5941158, 0.4962231, 0.6891587, 0.6216003, 0.2351496, 0.2201288, 
    0.3320474, 0.203185, 0.3021797, 0.5435779, 0.875765, 0.7273651, 1.251864, 
    0.9950132, 0.5095341, 0.4807606, 0.5004917, 0.2218755, 0.9272333, 
    0.3412112, 0.8966986, 0.6250736, 0.2526803, 0.5615672, 0.6932021, 
    0.5630955, 0.3327925, 0.239477, 0.3377306, 0.7845749, 0.9469273, 
    0.715499, 0.3157103, 0.1179704, 0.8387173, 0.2224763, 0.4719347, 
    0.5025061, 0.7269072, 0.6696218, 0.2286531, 0.2448571, 0.282111, 
    0.2615377, 0.2223855, 0.1434069, 0.1688031,
  0.6593438, 0.3609636, 0.2674334, 0.7208009, 0.2211715, 0.3771244, 0.502105, 
    0.78563, 0.3791666, 0.6154537, 0.1714588, 0.8821526, 0.1644452, 
    0.6376624, 0.8189439, 0.6955386, 0.2300579, 0.1458532, 0.2022019, 
    0.5415791, 0.2772168, 0.7236987, 0.2269711, 0.6120422, 0.3991513, 
    0.2252939, 0.8783276, 0.2224808, 0.2418258, 0.2090024, 0.1685721, 
    0.2237664, 0.3532139, 0.1439701, 0.6661603, 0.1875535, 0.4924571, 
    0.9841146, 0.1712926, 0.9878223, 0.3184504, 0.3175349, 0.458364, 
    0.8091118, 0.4263323, 0.3287061, 0.9641117, 0.2955255, 0.6129987, 
    0.7493274, 0.1465542, 0.2836272, 0.8138912, 0.1751759, 0.8053584, 
    0.2262039, 0.3357672, 0.4342431, 0.6833856, 0.7623785, 1.054256, 
    0.9113811, 0.6944475, 0.5373439, 0.3324913, 0.5390173, 0.250742, 
    0.3017584, 0.3172254, 0.6338109, 0.2760623, 0.3768659, 0.324406, 
    0.8443461, 0.5644274, 0.2881272, 0.3096578, 0.619137, 0.6527753, 
    0.4864714, 0.2781581, 0.9833164, 0.1467627, 0.6454289, 0.2878882, 
    0.817261, 0.5940058, 0.8498452, 0.3222598, 0.2337891, 0.1406264, 
    0.2607847, 0.1779588, 0.2798218, 0.2264215, 0.2744119,
  0.3055394, 0.2923887, 0.5920243, 0.3510437, 0.7482433, 0.3939995, 
    0.2687896, 0.553323, 0.2781042, 0.4202462, 0.8255653, 0.1815193, 
    0.2089593, 0.8083507, 0.2364269, 0.3107083, 0.9195414, 0.1531171, 
    0.198031, 0.3650708, 0.4963799, 0.7914947, 0.2362839, 0.1904638, 
    0.3813348, 0.5249822, 0.3827663, 0.5056133, 0.2191088, 0.2782821, 
    0.5364606, 0.2720293, 0.5261379, 0.1339067, 0.237537, 0.196823, 
    0.2179878, 0.3874499, 0.2989043, 0.2640974, 0.2123961, 0.5683975, 
    0.8370518, 0.5701421, 0.7762449, 0.7231753, 0.7561485, 0.7816435, 
    0.749617, 0.5105657, 0.2628373, 0.1899802, 0.8739544, 0.2404225, 
    0.3234132, 0.1244354, 0.2961805, 0.6494125, 0.7514091, 0.9981682, 
    1.132978, 0.5222794, 0.5794176, 0.3648824, 0.3596523, 0.5020914, 
    0.7645478, 0.9855402, 0.2705429, 0.8571758, 0.5636833, 0.8625976, 
    0.5463556, 0.832848, 0.4834849, 0.2178168, 0.3354498, 0.3885076, 
    0.5910681, 0.4060864, 0.2416416, 0.3232178, 0.4318793, 0.3390348, 
    0.6309202, 0.7157029, 0.7199245, 0.5076233, 0.9713045, 0.1567058, 
    0.2094672, 0.296649, 0.3212895, 0.3388297, 0.1872596, 0.2566147,
  0.444454, 0.7820367, 0.3064266, 0.3244969, 0.5235528, 0.5432233, 0.3553139, 
    0.6082892, 0.2675404, 0.1990476, 0.2439513, 0.1817257, 0.2853151, 
    0.823241, 0.2050045, 0.8546315, 0.3316197, 0.931179, 0.27967, 0.8770651, 
    0.5749466, 0.5448424, 0.2458876, 0.2694567, 0.8322615, 0.6623248, 
    0.747642, 0.3149025, 0.2847995, 0.2208068, 0.3111832, 0.3744749, 
    0.7674193, 0.3298192, 0.144244, 0.2095633, 0.3939396, 0.745603, 0.399391, 
    0.9490491, 0.4849875, 0.4606508, 0.3306073, 0.2158446, 0.3472773, 
    0.5323187, 0.5053442, 0.5432568, 0.3482898, 0.3217087, 0.1459292, 
    0.7416025, 0.8111308, 0.1594505, 0.2638705, 0.6749451, 0.836911, 
    0.5637347, 0.5239038, 0.7214295, 0.6195818, 0.392153, 0.4185706, 
    0.5075769, 0.192627, 0.1241125, 0.7334284, 0.3360943, 0.7594332, 
    0.6575118, 0.3842941, 0.9002581, 0.7779141, 0.812569, 0.4305702, 
    0.2334919, 0.2789024, 0.4420422, 0.530598, 0.3150181, 0.360597, 0.426633, 
    0.4628402, 0.7196789, 0.5608602, 0.7547588, 0.489637, 0.4729998, 
    0.3833358, 0.2931899, 0.2370045, 0.3119648, 0.4237458, 0.2278187, 
    0.1796433, 0.1323241,
  0.8491501, 0.6006591, 0.2254138, 0.7801049, 0.8244215, 0.558607, 0.5412297, 
    0.1992026, 0.8616919, 0.7105308, 0.417144, 0.1909727, 0.6804634, 
    0.7274687, 0.4305487, 0.9355896, 0.6633238, 0.9243693, 0.1222859, 
    0.2062387, 0.5457674, 0.9986019, 0.7826542, 0.7531931, 0.3431364, 
    0.1139358, 0.2618915, 0.1920516, 0.2145903, 0.2357506, 0.2740792, 
    0.5600311, 0.7589592, 0.8606415, 0.915633, 0.1969787, 0.3631368, 
    0.6161781, 0.2787137, 0.9348773, 0.336744, 0.621555, 0.9225765, 
    0.3690377, 0.4155008, 0.5254639, 0.2412468, 0.2071874, 0.2439197, 
    0.4940676, 0.4828147, 0.4342853, 0.4137139, 0.8020678, 0.6085526, 
    0.7929617, 0.9532921, 0.5282161, 0.5780501, 0.5261132, 0.783304, 
    0.4321966, 0.4456051, 0.4903353, 0.8211594, 0.6384828, 0.2323455, 
    0.4458759, 0.9174932, 0.4980997, 0.6074433, 0.7582713, 0.8228168, 
    0.6124404, 0.6034449, 0.5235595, 0.3870348, 0.3784181, 0.4548996, 
    0.540296, 0.7773914, 0.7053837, 0.4292297, 0.612976, 0.5201478, 
    0.4238658, 0.6445412, 0.3252737, 0.3647941, 0.1613467, 0.2405015, 
    0.3335114, 0.3071654, 0.3259597, 0.4628202, 0.1670586,
  0.663556, 0.6732333, 0.1863649, 0.6056557, 0.4877072, 0.42026, 0.3057786, 
    0.4889986, 0.5255104, 0.9034796, 0.231222, 0.2384451, 0.2327916, 
    0.5214932, 0.7483705, 0.8207703, 0.5488306, 0.8845263, 0.432458, 0.8653, 
    0.2752009, 0.6616606, 0.2609529, 0.4626007, 0.7971273, 0.2366795, 
    0.1483282, 0.1714887, 0.3035242, 0.2769368, 0.9368467, 0.5783767, 
    0.3526831, 0.7464561, 0.8298263, 0.2976183, 0.2062079, 0.3416952, 
    0.5108322, 0.2983678, 0.5105064, 0.5971901, 0.3414758, 0.4461374, 
    0.6933995, 0.5367584, 0.5432771, 0.6129616, 0.4668052, 0.7196918, 
    0.8732188, 0.6541534, 0.5996124, 0.2179756, 0.85923, 0.4586002, 
    0.9400957, 0.4443735, 0.2959612, 0.8897257, 0.4961368, 0.3911729, 
    0.7337782, 0.3838522, 0.2833546, 0.2278309, 0.3855826, 0.534655, 
    0.8938532, 0.2890951, 0.1388913, 0.1946098, 0.4333963, 0.6614031, 
    0.4874207, 0.48159, 0.3502133, 0.3501068, 0.5339236, 0.7125043, 
    0.7735588, 0.5690976, 0.4292995, 0.650019, 0.4812855, 0.3700157, 
    0.3301862, 0.4230283, 0.3129591, 0.1626379, 0.09073837, 0.3392093, 
    0.5095114, 0.5757693, 0.6860257, 0.5187959,
  0.5705903, 0.4820425, 0.4467522, 0.3837257, 0.3589422, 0.2269406, 
    0.3691883, 0.3211596, 0.9802056, 0.4748353, 0.2449672, 0.25946, 
    0.8244318, 0.6646013, 0.8296453, 0.4414392, 0.5037096, 0.7456715, 
    0.6025747, 0.4854253, 0.1992539, 0.585939, 0.3550005, 0.5174885, 
    0.9229558, 0.6628724, 0.6770101, 0.2924789, 0.352128, 0.1989041, 
    0.9079929, 0.3879872, 0.6676182, 0.4728896, 0.2988791, 0.1401567, 
    0.1248084, 0.8174673, 0.3541858, 0.2688991, 0.3318263, 0.3120928, 
    0.4395972, 0.3852765, 0.694636, 0.4572604, 0.6873885, 0.6204996, 
    0.2370412, 0.321958, 0.8780817, 0.2731156, 0.2258738, 0.3088748, 
    0.7131113, 0.4756933, 0.4459488, 0.3359571, 0.7280603, 0.5205888, 
    0.5004314, 0.4702863, 0.8700247, 0.3669756, 0.2704104, 0.3901683, 
    0.3120538, 0.3529272, 0.7064658, 0.1157412, 0.1874142, 0.3531048, 
    0.7482743, 0.6253453, 0.5600945, 0.3267074, 0.2621759, 0.2653536, 
    0.4670306, 0.878021, 0.4656478, 0.5430589, 0.3221894, 0.5362661, 
    0.350185, 0.3480993, 0.4326323, 0.4660952, 0.4469193, 0.1495365, 
    0.2237365, 0.4096938, 0.4775677, 0.9781163, 0.4854324, 0.4679533 ;

 CldBase =
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888 ;

 CldThick =
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888 ;

 CldTop =
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888 ;

 Emis =
  8713, 8824, 8958, 8960, 8962, 8964, 8966, 8967, 8968, 8971, 8971, 8971, 
    8971, 8971, 8971, 8994, 9086, 9086, 9086, 9086, 9086, 9086,
  8757, 8863, 8964, 8965, 8966, 8966, 8967, 8968, 8968, 8969, 8969, 8969, 
    8969, 8969, 8969, 8977, 9014, 9014, 9014, 9014, 9014, 9014,
  8913, 9015, 9093, 9092, 9091, 9090, 9091, 9090, 9090, 9088, 9088, 9088, 
    9088, 9088, 9088, 9086, 9048, 9048, 9048, 9048, 9048, 9048,
  8942, 9040, 9121, 9122, 9123, 9123, 9124, 9124, 9125, 9126, 9126, 9126, 
    9126, 9126, 9126, 9114, 9162, 9162, 9162, 9162, 9162, 9162,
  8876, 8975, 9002, 9004, 9005, 9006, 9008, 9009, 9010, 9012, 9012, 9012, 
    9012, 9012, 9012, 9037, 9097, 9097, 9097, 9097, 9097, 9097,
  8860, 8961, 8972, 8975, 8978, 8979, 8982, 8983, 8984, 8988, 8988, 8988, 
    8988, 8988, 8988, 9038, 9121, 9121, 9121, 9121, 9122, 9121,
  8912, 9013, 9017, 9018, 9019, 9019, 9021, 9021, 9022, 9023, 9023, 9023, 
    9023, 9023, 9023, 9066, 9079, 9079, 9079, 9079, 9079, 9079,
  8864, 8969, 8914, 8913, 8913, 8912, 8913, 8913, 8912, 8911, 8911, 8911, 
    8911, 8911, 8911, 8990, 8889, 8889, 8889, 8889, 8889, 8889,
  8949, 9050, 8977, 8977, 8977, 8977, 8977, 8977, 8977, 8977, 8977, 8977, 
    8977, 8977, 8977, 9053, 8987, 8987, 8987, 8987, 8987, 8987,
  8964, 9052, 8864, 8857, 8851, 8847, 8844, 8841, 8838, 8830, 8830, 8830, 
    8830, 8830, 8830, 8864, 8549, 8549, 8549, 8549, 8549, 8549,
  8999, 9098, 8993, 8993, 8993, 8993, 8994, 8993, 8993, 8993, 8993, 8993, 
    8993, 8993, 8993, 9073, 8992, 8992, 8992, 8992, 8992, 8992,
  8993, 9093, 8975, 8976, 8977, 8978, 8980, 8980, 8981, 8983, 8983, 8983, 
    8983, 8983, 8983, 9090, 9053, 9053, 9053, 9053, 9053, 9053,
  9078, 9172, 9007, 9008, 9008, 9009, 9010, 9010, 9011, 9012, 9012, 9012, 
    9012, 9012, 9012, 9113, 9052, 9052, 9052, 9052, 9052, 9052,
  8995, 9095, 9042, 9043, 9043, 9044, 9045, 9045, 9046, 9047, 9047, 9047, 
    9047, 9047, 9047, 9119, 9090, 9090, 9090, 9090, 9090, 9090,
  8766, 8874, 8741, 8738, 8737, 8735, 8735, 8734, 8733, 8731, 8731, 8731, 
    8731, 8731, 8731, 8846, 8651, 8651, 8651, 8651, 8651, 8651,
  9161, 9234, 8953, 8943, 8936, 8931, 8926, 8923, 8919, 8908, 8908, 8908, 
    8908, 8908, 8908, 8913, 8549, 8549, 8549, 8549, 8549, 8549,
  9128, 9206, 8866, 8858, 8853, 8849, 8846, 8843, 8841, 8832, 8832, 8832, 
    8832, 8832, 8832, 8904, 8560, 8560, 8560, 8560, 8560, 8560,
  9062, 9150, 8875, 8868, 8862, 8858, 8855, 8852, 8849, 8840, 8840, 8840, 
    8840, 8840, 8840, 8917, 8559, 8559, 8559, 8559, 8559, 8559,
  9092, 9187, 8931, 8931, 8931, 8931, 8932, 8932, 8932, 8932, 8932, 8932, 
    8932, 8932, 8932, 9080, 8939, 8939, 8939, 8939, 8939, 8939,
  9107, 9204, 8959, 8962, 8963, 8964, 8966, 8967, 8968, 8970, 8970, 8970, 
    8970, 8970, 8970, 9133, 9060, 9060, 9060, 9060, 9060, 9060,
  9002, 9095, 8769, 8767, 8765, 8764, 8764, 8763, 8762, 8759, 8759, 8759, 
    8759, 8759, 8759, 8920, 8683, 8683, 8683, 8683, 8683, 8683,
  9054, 9150, 8816, 8814, 8813, 8813, 8813, 8813, 8812, 8811, 8811, 8811, 
    8811, 8811, 8811, 8996, 8771, 8771, 8771, 8771, 8771, 8771,
  9056, 9156, 8744, 8743, 8743, 8743, 8744, 8744, 8744, 8743, 8743, 8743, 
    8743, 8743, 8743, 8989, 8741, 8741, 8741, 8741, 8741, 8741,
  9079, 9176, 8766, 8764, 8763, 8762, 8762, 8762, 8761, 8759, 8759, 8759, 
    8759, 8759, 8759, 8985, 8706, 8706, 8706, 8706, 8706, 8706,
  9082, 9177, 8787, 8787, 8786, 8786, 8786, 8786, 8786, 8785, 8785, 8785, 
    8785, 8785, 8785, 8999, 8770, 8770, 8770, 8770, 8770, 8770,
  9046, 9141, 8763, 8762, 8761, 8761, 8762, 8762, 8761, 8761, 8761, 8761, 
    8761, 8761, 8761, 8970, 8746, 8746, 8746, 8746, 8746, 8746,
  9172, 9259, 8911, 8909, 8908, 8907, 8906, 8906, 8905, 8902, 8902, 8902, 
    8902, 8902, 8902, 9054, 8831, 8831, 8831, 8831, 8831, 8831,
  9196, 9282, 8886, 8883, 8882, 8880, 8880, 8879, 8878, 8875, 8875, 8875, 
    8875, 8875, 8875, 9042, 8787, 8787, 8787, 8787, 8787, 8787,
  9252, 9337, 8921, 8919, 8917, 8916, 8915, 8914, 8913, 8911, 8911, 8911, 
    8911, 8911, 8911, 9087, 8829, 8829, 8829, 8829, 8829, 8829,
  9185, 9273, 8883, 8881, 8880, 8879, 8878, 8878, 8877, 8875, 8875, 8875, 
    8875, 8875, 8875, 9055, 8808, 8808, 8808, 8808, 8808, 8808,
  9128, 9220, 8827, 8826, 8825, 8825, 8825, 8825, 8824, 8823, 8823, 8823, 
    8823, 8823, 8823, 9026, 8793, 8793, 8793, 8793, 8793, 8793,
  9053, 9151, 8756, 8756, 8755, 8755, 8756, 8756, 8756, 8756, 8756, 8756, 
    8756, 8756, 8756, 8988, 8755, 8755, 8755, 8755, 8755, 8755,
  9091, 9182, 8785, 8785, 8784, 8784, 8784, 8784, 8784, 8783, 8783, 8783, 
    8783, 8783, 8783, 8981, 8763, 8763, 8763, 8763, 8763, 8763,
  8507, 8632, 8227, 8231, 8234, 8236, 8239, 8240, 8242, 8246, 8246, 8246, 
    8246, 8246, 8246, 8609, 8398, 8398, 8398, 8398, 8398, 8398,
  8270, 8406, 8123, 8128, 8132, 8135, 8138, 8140, 8142, 8148, 8148, 8148, 
    8148, 8148, 8148, 8496, 8354, 8354, 8354, 8354, 8354, 8354,
  8331, 8464, 8212, 8217, 8220, 8223, 8226, 8228, 8229, 8235, 8235, 8235, 
    8235, 8235, 8235, 8551, 8418, 8418, 8418, 8418, 8418, 8418,
  8238, 8379, 8044, 8050, 8055, 8058, 8063, 8065, 8067, 8075, 8075, 8075, 
    8075, 8075, 8075, 8481, 8329, 8329, 8329, 8329, 8329, 8329,
  8563, 8684, 8439, 8441, 8443, 8444, 8447, 8448, 8449, 8451, 8451, 8451, 
    8451, 8451, 8451, 8707, 8558, 8558, 8558, 8558, 8558, 8558,
  8391, 8520, 8208, 8211, 8214, 8215, 8218, 8219, 8220, 8223, 8223, 8223, 
    8223, 8223, 8223, 8550, 8346, 8346, 8346, 8346, 8346, 8346,
  8488, 8608, 8456, 8455, 8454, 8453, 8453, 8453, 8452, 8451, 8451, 8451, 
    8451, 8451, 8451, 8630, 8410, 8410, 8410, 8410, 8410, 8410,
  8339, 8466, 8287, 8288, 8289, 8290, 8291, 8292, 8292, 8293, 8293, 8293, 
    8293, 8293, 8293, 8526, 8345, 8345, 8345, 8345, 8345, 8345,
  8386, 8522, 8293, 8297, 8300, 8302, 8305, 8307, 8308, 8312, 8312, 8312, 
    8312, 8312, 8312, 8633, 8471, 8471, 8471, 8471, 8471, 8471,
  8371, 8510, 8134, 8140, 8144, 8147, 8151, 8153, 8155, 8162, 8162, 8162, 
    8162, 8162, 8162, 8578, 8390, 8390, 8390, 8390, 8390, 8390,
  8459, 8594, 8218, 8221, 8224, 8226, 8229, 8230, 8231, 8235, 8235, 8235, 
    8235, 8235, 8235, 8625, 8380, 8380, 8380, 8380, 8380, 8380,
  8324, 8464, 8113, 8116, 8118, 8120, 8122, 8123, 8124, 8128, 8128, 8128, 
    8128, 8128, 8128, 8515, 8251, 8251, 8251, 8251, 8251, 8251,
  8384, 8519, 8225, 8226, 8227, 8228, 8229, 8230, 8230, 8232, 8232, 8232, 
    8232, 8232, 8232, 8563, 8294, 8294, 8294, 8294, 8294, 8294,
  8502, 8641, 8412, 8416, 8418, 8420, 8423, 8424, 8426, 8430, 8430, 8430, 
    8430, 8430, 8430, 8765, 8577, 8577, 8577, 8577, 8577, 8577,
  8449, 8580, 8252, 8252, 8252, 8252, 8253, 8253, 8253, 8252, 8252, 8252, 
    8252, 8252, 8252, 8575, 8260, 8260, 8260, 8260, 8260, 8260,
  8473, 8598, 8218, 8216, 8214, 8213, 8213, 8213, 8212, 8209, 8209, 8209, 
    8209, 8209, 8209, 8520, 8144, 8144, 8144, 8144, 8144, 8144,
  8288, 8422, 8268, 8272, 8275, 8278, 8281, 8283, 8284, 8289, 8289, 8289, 
    8289, 8289, 8289, 8556, 8468, 8468, 8468, 8468, 8468, 8468,
  8605, 8746, 8442, 8445, 8448, 8450, 8453, 8454, 8455, 8459, 8459, 8459, 
    8459, 8459, 8459, 8843, 8607, 8607, 8607, 8607, 8607, 8607,
  8530, 8664, 8364, 8369, 8372, 8374, 8378, 8379, 8381, 8386, 8386, 8386, 
    8386, 8386, 8386, 8738, 8562, 8562, 8562, 8562, 8562, 8562,
  8444, 8581, 8345, 8349, 8353, 8355, 8358, 8360, 8362, 8367, 8367, 8367, 
    8367, 8367, 8367, 8699, 8547, 8547, 8547, 8547, 8547, 8547,
  8349, 8485, 8345, 8349, 8352, 8354, 8357, 8359, 8360, 8365, 8365, 8365, 
    8365, 8365, 8365, 8634, 8529, 8529, 8529, 8529, 8529, 8529,
  8254, 8395, 8180, 8184, 8187, 8189, 8193, 8194, 8196, 8201, 8201, 8201, 
    8201, 8201, 8201, 8530, 8377, 8377, 8377, 8377, 8377, 8377,
  8157, 8311, 8000, 8013, 8023, 8030, 8038, 8043, 8048, 8063, 8063, 8063, 
    8063, 8063, 8063, 8547, 8578, 8578, 8578, 8578, 8578, 8578,
  7825, 7994, 7691, 7716, 7734, 7747, 7761, 7770, 7779, 7807, 7807, 7807, 
    7807, 7807, 7807, 8413, 8753, 8753, 8753, 8753, 8753, 8753,
  7385, 7574, 7480, 7511, 7532, 7549, 7566, 7577, 7588, 7622, 7622, 7622, 
    7622, 7622, 7622, 8230, 8785, 8785, 8785, 8785, 8785, 8785,
  6949, 7159, 6978, 7006, 7026, 7041, 7058, 7068, 7078, 7110, 7110, 7110, 
    7110, 7110, 7110, 7829, 8188, 8188, 8188, 8188, 8188, 8188,
  6567, 6745, 6372, 6415, 6445, 6467, 6489, 6504, 6519, 6566, 6566, 6566, 
    6566, 6566, 6566, 7514, 8150, 8150, 8150, 8150, 8150, 8150,
  5966, 6135, 5565, 5614, 5649, 5674, 5700, 5716, 5734, 5788, 5788, 5788, 
    5788, 5788, 5788, 6996, 7608, 7608, 7608, 7608, 7608, 7608,
  5353, 5624, 5560, 5596, 5621, 5641, 5660, 5672, 5686, 5728, 5728, 5728, 
    5728, 5728, 5728, 6947, 7250, 7404, 7404, 7404, 7404, 7404,
  5086, 5376, 5476, 5514, 5542, 5563, 5583, 5596, 5611, 5655, 5655, 5655, 
    5655, 5655, 5655, 6781, 7237, 7393, 7393, 7393, 7393, 7393,
  5208, 5483, 5513, 5550, 5576, 5596, 5615, 5628, 5642, 5684, 5684, 5684, 
    5684, 5684, 5684, 6827, 7220, 7374, 7374, 7374, 7374, 7374,
  5557, 5816, 5802, 5836, 5860, 5878, 5896, 5907, 5921, 5960, 5960, 5960, 
    5960, 5960, 5960, 7060, 7379, 7525, 7525, 7525, 7525, 7525,
  5940, 6181, 6207, 6237, 6259, 6275, 6291, 6302, 6314, 6349, 6349, 6349, 
    6349, 6349, 6349, 7299, 7614, 7748, 7748, 7748, 7748, 7748,
  6276, 6515, 6608, 6637, 6657, 6673, 6688, 6697, 6709, 6741, 6741, 6741, 
    6741, 6741, 6741, 7563, 7890, 8013, 8013, 8013, 8013, 8013,
  6600, 6823, 6888, 6914, 6933, 6946, 6960, 6969, 6979, 7008, 7008, 7008, 
    7008, 7008, 7008, 7772, 8042, 8157, 8157, 8157, 8157, 8157,
  6837, 7056, 7007, 7032, 7050, 7063, 7076, 7084, 7094, 7122, 7122, 7122, 
    7122, 7122, 7122, 7967, 8116, 8229, 8229, 8229, 8229, 8229,
  6949, 7158, 7065, 7088, 7105, 7117, 7130, 7137, 7147, 7173, 7173, 7173, 
    7173, 7173, 7173, 8025, 8132, 8243, 8243, 8243, 8243, 8243,
  6948, 7135, 6873, 6895, 6911, 6923, 6934, 6941, 6950, 6976, 6976, 6976, 
    6976, 6976, 6976, 7961, 7947, 8063, 8063, 8063, 8063, 8063,
  6899, 7090, 6869, 6891, 6908, 6920, 6931, 6939, 6948, 6974, 6974, 6974, 
    6974, 6974, 6974, 7933, 7956, 8073, 8073, 8073, 8073, 8073,
  6793, 7002, 6908, 6932, 6950, 6963, 6975, 6984, 6993, 7021, 7021, 7021, 
    7021, 7021, 7021, 7900, 8027, 8143, 8143, 8143, 8143, 8143,
  6626, 6863, 6819, 6846, 6866, 6881, 6895, 6904, 6915, 6946, 6946, 6946, 
    6946, 6946, 6946, 7865, 8035, 8153, 8153, 8153, 8153, 8153,
  6420, 6654, 6614, 6641, 6661, 6676, 6691, 6700, 6711, 6743, 6743, 6743, 
    6743, 6743, 6743, 7681, 7879, 8002, 8002, 8002, 8002, 8002,
  6143, 6393, 6332, 6363, 6384, 6401, 6417, 6428, 6440, 6475, 6475, 6475, 
    6475, 6475, 6475, 7521, 7730, 7862, 7862, 7862, 7862, 7862,
  5797, 6067, 6006, 6040, 6065, 6083, 6101, 6113, 6126, 6165, 6165, 6165, 
    6165, 6165, 6165, 7312, 7555, 7697, 7697, 7697, 7697, 7697,
  5441, 5718, 5568, 5605, 5631, 5650, 5669, 5682, 5696, 5738, 5738, 5738, 
    5738, 5738, 5738, 7058, 7271, 7426, 7426, 7426, 7426, 7426,
  5149, 5432, 5328, 5366, 5394, 5414, 5434, 5448, 5462, 5507, 5507, 5507, 
    5507, 5507, 5507, 6834, 7118, 7279, 7279, 7279, 7279, 7279,
  4969, 5249, 5232, 5270, 5297, 5318, 5338, 5352, 5367, 5411, 5411, 5411, 
    5411, 5411, 5411, 6657, 7038, 7200, 7200, 7200, 7200, 7200,
  5012, 5297, 5237, 5276, 5304, 5325, 5345, 5359, 5373, 5418, 5418, 5418, 
    5418, 5418, 5418, 6720, 7057, 7220, 7220, 7220, 7220, 7220,
  5294, 5596, 5588, 5627, 5655, 5676, 5696, 5710, 5725, 5770, 5770, 5770, 
    5770, 5770, 5770, 7021, 7353, 7509, 7509, 7509, 7509, 7509,
  5961, 6228, 6209, 6242, 6265, 6283, 6300, 6312, 6324, 6362, 6362, 6362, 
    6362, 6362, 6362, 7431, 7689, 7825, 7825, 7825, 7825, 7825,
  6620, 6830, 6957, 6981, 6999, 7012, 7025, 7033, 7042, 7070, 7070, 7070, 
    7070, 7070, 7070, 7724, 8052, 8164, 8164, 8164, 8164, 8164,
  7188, 7374, 7494, 7513, 7528, 7538, 7548, 7555, 7563, 7585, 7585, 7585, 
    7585, 7585, 7585, 8099, 8363, 8458, 8458, 8458, 8458, 8458,
  7633, 7776, 7777, 7790, 7800, 7808, 7815, 7819, 7826, 7841, 7841, 7841, 
    7841, 7841, 7841, 8307, 8443, 8529, 8529, 8529, 8529, 8529,
  7941, 8185, 8197, 8202, 8206, 8208, 8211, 8212, 8214, 8220, 8220, 8220, 
    8220, 8220, 8220, 8546, 8405, 8405, 8405, 8405, 8405, 8405,
  7958, 8174, 8145, 8149, 8152, 8154, 8156, 8157, 8159, 8163, 8163, 8163, 
    8163, 8163, 8163, 8434, 8310, 8310, 8310, 8310, 8310, 8310,
  7946, 8063, 8066, 8075, 8083, 8088, 8094, 8097, 8101, 8113, 8113, 8113, 
    8113, 8113, 8113, 8459, 8573, 8649, 8649, 8649, 8649, 8649,
  7781, 7944, 8122, 8131, 8137, 8142, 8147, 8150, 8153, 8163, 8163, 8163, 
    8163, 8163, 8163, 8399, 8503, 8503, 8503, 8503, 8503, 8503,
  7811, 7972, 8153, 8162, 8168, 8173, 8179, 8182, 8185, 8195, 8195, 8195, 
    8195, 8195, 8195, 8424, 8545, 8545, 8545, 8545, 8545, 8545,
  7989, 8270, 8475, 8467, 8461, 8456, 8452, 8448, 8445, 8435, 8435, 8435, 
    8435, 8435, 8435, 8515, 8107, 8107, 8107, 8107, 8107, 8107,
  7838, 8129, 8444, 8431, 8423, 8416, 8409, 8405, 8400, 8386, 8386, 8386, 
    8386, 8386, 8386, 8334, 7911, 7911, 7911, 7911, 7911, 7911,
  7533, 7790, 8076, 8066, 8060, 8054, 8049, 8045, 8041, 8030, 8030, 8030, 
    8030, 8030, 8030, 7922, 7648, 7648, 7648, 7648, 7648, 7648,
  7130, 7473, 7988, 7978, 7971, 7966, 7961, 7956, 7953, 7941, 7941, 7941, 
    7941, 7941, 7941, 7856, 7559, 7559, 7559, 7559, 7559, 7559,
  6925, 7370, 8115, 8102, 8093, 8085, 8078, 8073, 8068, 8053, 8053, 8053, 
    8053, 8053, 8053, 8004, 7549, 7549, 7549, 7549, 7549, 7549,
  8727, 8840, 8997, 8999, 9001, 9002, 9004, 9005, 9005, 9008, 9008, 9008, 
    9008, 9008, 9008, 9025, 9094, 9094, 9094, 9094, 9094, 9094,
  8789, 8897, 9022, 9023, 9024, 9025, 9027, 9027, 9028, 9029, 9029, 9029, 
    9029, 9029, 9029, 9040, 9091, 9091, 9091, 9091, 9091, 9091,
  8903, 9010, 9073, 9067, 9063, 9060, 9058, 9056, 9054, 9047, 9047, 9047, 
    9047, 9047, 9047, 9045, 8844, 8844, 8844, 8844, 8844, 8844,
  8969, 9068, 9178, 9176, 9175, 9174, 9174, 9173, 9172, 9170, 9170, 9170, 
    9170, 9170, 9170, 9133, 9105, 9105, 9105, 9105, 9105, 9105,
  8974, 9076, 9141, 9141, 9142, 9142, 9143, 9143, 9144, 9144, 9144, 9144, 
    9144, 9144, 9144, 9161, 9178, 9178, 9178, 9178, 9178, 9178,
  8887, 8991, 9020, 9022, 9023, 9024, 9026, 9026, 9027, 9029, 9029, 9029, 
    9029, 9029, 9029, 9076, 9104, 9104, 9104, 9104, 9104, 9104,
  9005, 9106, 9035, 9035, 9035, 9034, 9035, 9035, 9035, 9035, 9035, 9035, 
    9035, 9035, 9035, 9109, 9034, 9034, 9034, 9034, 9034, 9034,
  9001, 9096, 9010, 9007, 9004, 9002, 9001, 9000, 8999, 8995, 8995, 8995, 
    8995, 8995, 8995, 9032, 8871, 8871, 8871, 8871, 8871, 8871,
  9153, 9228, 9128, 9116, 9107, 9101, 9095, 9091, 9086, 9073, 9073, 9073, 
    9073, 9073, 9073, 8981, 8628, 8628, 8628, 8628, 8628, 8628,
  8980, 9080, 8990, 8990, 8991, 8991, 8992, 8992, 8992, 8993, 8993, 8993, 
    8993, 8993, 8993, 9080, 9021, 9021, 9021, 9021, 9021, 9021,
  9014, 9112, 8955, 8957, 8957, 8958, 8960, 8960, 8960, 8962, 8962, 8962, 
    8962, 8962, 8962, 9075, 9014, 9014, 9014, 9014, 9014, 9014,
  9021, 9119, 8934, 8935, 8936, 8937, 8939, 8939, 8940, 8942, 8942, 8942, 
    8942, 8942, 8942, 9073, 9009, 9009, 9009, 9009, 9009, 9009,
  8944, 9047, 8961, 8963, 8964, 8965, 8967, 8967, 8968, 8970, 8970, 8970, 
    8970, 8970, 8970, 9071, 9048, 9048, 9048, 9048, 9048, 9048,
  9091, 9181, 8984, 8983, 8982, 8981, 8982, 8981, 8981, 8980, 8980, 8980, 
    8980, 8980, 8980, 9074, 8949, 8949, 8949, 8949, 8949, 8949,
  8808, 8913, 8685, 8683, 8681, 8680, 8679, 8678, 8678, 8675, 8675, 8675, 
    8675, 8675, 8675, 8831, 8593, 8593, 8593, 8593, 8593, 8593,
  8823, 8931, 8603, 8602, 8601, 8600, 8601, 8600, 8600, 8598, 8598, 8598, 
    8598, 8598, 8598, 8824, 8558, 8558, 8558, 8558, 8558, 8558,
  8931, 9037, 8679, 8679, 8679, 8678, 8679, 8679, 8679, 8678, 8678, 8678, 
    8678, 8678, 8678, 8920, 8673, 8673, 8673, 8673, 8673, 8673,
  8989, 9083, 8712, 8708, 8706, 8704, 8703, 8702, 8700, 8696, 8696, 8696, 
    8696, 8696, 8696, 8878, 8574, 8574, 8574, 8574, 8574, 8574,
  9005, 9096, 8769, 8765, 8763, 8761, 8761, 8760, 8758, 8755, 8755, 8755, 
    8755, 8755, 8755, 8899, 8645, 8645, 8645, 8645, 8645, 8645,
  9072, 9162, 8881, 8873, 8866, 8862, 8858, 8855, 8852, 8842, 8842, 8842, 
    8842, 8842, 8842, 8927, 8523, 8523, 8523, 8523, 8523, 8523,
  9012, 9104, 8836, 8833, 8832, 8830, 8830, 8829, 8828, 8826, 8826, 8826, 
    8826, 8826, 8826, 8951, 8748, 8748, 8748, 8748, 8748, 8748,
  9068, 9160, 8846, 8842, 8839, 8837, 8836, 8835, 8833, 8829, 8829, 8829, 
    8829, 8829, 8829, 8967, 8689, 8689, 8689, 8689, 8689, 8689,
  9029, 9126, 8757, 8754, 8752, 8751, 8751, 8750, 8749, 8746, 8746, 8746, 
    8746, 8746, 8746, 8940, 8658, 8658, 8658, 8658, 8658, 8658,
  9124, 9218, 8825, 8822, 8820, 8819, 8819, 8818, 8817, 8814, 8814, 8814, 
    8814, 8814, 8814, 9012, 8725, 8725, 8725, 8725, 8725, 8725,
  9024, 9124, 8700, 8701, 8701, 8701, 8702, 8702, 8702, 8703, 8703, 8703, 
    8703, 8703, 8703, 8962, 8724, 8724, 8724, 8724, 8724, 8724,
  9016, 9115, 8738, 8738, 8738, 8738, 8739, 8739, 8739, 8738, 8738, 8738, 
    8738, 8738, 8738, 8964, 8746, 8746, 8746, 8746, 8746, 8746,
  9103, 9196, 8810, 8809, 8808, 8808, 8808, 8808, 8807, 8806, 8806, 8806, 
    8806, 8806, 8806, 9010, 8779, 8779, 8779, 8779, 8779, 8779,
  9242, 9327, 8941, 8939, 8938, 8936, 8936, 8936, 8935, 8932, 8932, 8932, 
    8932, 8932, 8932, 9093, 8862, 8862, 8862, 8862, 8862, 8862,
  9295, 9379, 8976, 8972, 8970, 8968, 8968, 8966, 8965, 8961, 8961, 8961, 
    8961, 8961, 8961, 9125, 8848, 8848, 8848, 8848, 8848, 8848,
  9175, 9264, 8870, 8867, 8865, 8863, 8862, 8861, 8860, 8857, 8857, 8857, 
    8857, 8857, 8857, 9037, 8748, 8748, 8748, 8748, 8748, 8748,
  9031, 9130, 8715, 8715, 8715, 8715, 8716, 8716, 8716, 8716, 8716, 8716, 
    8716, 8716, 8716, 8962, 8727, 8727, 8727, 8727, 8727, 8727,
  8980, 9083, 8644, 8645, 8645, 8646, 8647, 8647, 8648, 8649, 8649, 8649, 
    8649, 8649, 8649, 8927, 8687, 8687, 8687, 8687, 8687, 8687,
  8969, 9069, 8689, 8689, 8689, 8689, 8690, 8690, 8690, 8690, 8690, 8690, 
    8690, 8690, 8690, 8923, 8708, 8708, 8708, 8708, 8708, 8708,
  8745, 8856, 8544, 8546, 8547, 8548, 8549, 8550, 8550, 8552, 8552, 8552, 
    8552, 8552, 8552, 8801, 8620, 8620, 8620, 8620, 8620, 8620,
  8643, 8759, 8501, 8503, 8505, 8506, 8508, 8509, 8510, 8512, 8512, 8512, 
    8512, 8512, 8512, 8757, 8608, 8608, 8608, 8608, 8608, 8608,
  8407, 8538, 8317, 8320, 8323, 8324, 8327, 8329, 8330, 8334, 8334, 8334, 
    8334, 8334, 8334, 8624, 8476, 8476, 8476, 8476, 8476, 8476,
  8339, 8474, 8239, 8242, 8245, 8247, 8250, 8252, 8253, 8257, 8257, 8257, 
    8257, 8257, 8257, 8569, 8413, 8413, 8413, 8413, 8413, 8413,
  8294, 8429, 8153, 8158, 8161, 8163, 8167, 8168, 8170, 8175, 8175, 8175, 
    8175, 8175, 8175, 8513, 8358, 8358, 8358, 8358, 8358, 8358,
  8434, 8562, 8328, 8331, 8333, 8334, 8337, 8338, 8339, 8342, 8342, 8342, 
    8342, 8342, 8342, 8624, 8462, 8462, 8462, 8462, 8462, 8462,
  8317, 8446, 8201, 8203, 8205, 8206, 8208, 8209, 8210, 8213, 8213, 8213, 
    8213, 8213, 8213, 8498, 8311, 8311, 8311, 8311, 8311, 8311,
  8258, 8394, 8202, 8207, 8210, 8213, 8216, 8218, 8219, 8224, 8224, 8224, 
    8224, 8224, 8224, 8522, 8404, 8404, 8404, 8404, 8404, 8404,
  8508, 8636, 8273, 8275, 8276, 8277, 8280, 8280, 8281, 8284, 8284, 8284, 
    8284, 8284, 8284, 8631, 8376, 8376, 8376, 8376, 8376, 8376,
  8528, 8659, 8223, 8228, 8231, 8233, 8236, 8238, 8239, 8244, 8244, 8244, 
    8244, 8244, 8244, 8650, 8418, 8418, 8418, 8418, 8418, 8418,
  8457, 8591, 8155, 8159, 8162, 8164, 8167, 8168, 8170, 8174, 8174, 8174, 
    8174, 8174, 8174, 8593, 8335, 8335, 8335, 8335, 8335, 8335,
  8499, 8630, 8259, 8262, 8264, 8266, 8268, 8270, 8270, 8274, 8274, 8274, 
    8274, 8274, 8274, 8641, 8394, 8394, 8394, 8394, 8394, 8394,
  8499, 8629, 8338, 8338, 8338, 8339, 8340, 8340, 8340, 8341, 8341, 8341, 
    8341, 8341, 8341, 8647, 8370, 8370, 8370, 8370, 8370, 8370,
  8499, 8625, 8456, 8455, 8454, 8454, 8454, 8454, 8453, 8452, 8452, 8452, 
    8452, 8452, 8452, 8669, 8419, 8419, 8419, 8419, 8419, 8419,
  8479, 8607, 8414, 8415, 8416, 8416, 8418, 8418, 8419, 8420, 8420, 8420, 
    8420, 8420, 8420, 8672, 8470, 8470, 8470, 8470, 8470, 8470,
  8579, 8708, 8314, 8318, 8321, 8323, 8326, 8328, 8329, 8333, 8333, 8333, 
    8333, 8333, 8333, 8711, 8488, 8488, 8488, 8488, 8488, 8488,
  8614, 8742, 8346, 8352, 8356, 8359, 8363, 8365, 8367, 8374, 8374, 8374, 
    8374, 8374, 8374, 8763, 8598, 8598, 8598, 8598, 8598, 8598,
  8479, 8607, 8235, 8240, 8243, 8245, 8248, 8250, 8252, 8257, 8257, 8257, 
    8257, 8257, 8257, 8617, 8433, 8433, 8433, 8433, 8433, 8433,
  8474, 8602, 8264, 8267, 8270, 8272, 8275, 8276, 8277, 8281, 8281, 8281, 
    8281, 8281, 8281, 8616, 8426, 8426, 8426, 8426, 8425, 8425,
  8502, 8628, 8346, 8350, 8353, 8354, 8357, 8359, 8360, 8364, 8364, 8364, 
    8364, 8364, 8364, 8663, 8512, 8512, 8512, 8512, 8512, 8512,
  8448, 8585, 8309, 8314, 8317, 8319, 8323, 8324, 8326, 8331, 8331, 8331, 
    8331, 8331, 8331, 8687, 8516, 8516, 8516, 8516, 8516, 8516,
  8363, 8505, 8265, 8270, 8273, 8275, 8278, 8280, 8281, 8286, 8286, 8286, 
    8286, 8286, 8286, 8635, 8458, 8458, 8458, 8458, 8458, 8458,
  8238, 8381, 8049, 8056, 8060, 8064, 8069, 8071, 8073, 8081, 8081, 8081, 
    8081, 8081, 8081, 8492, 8343, 8343, 8343, 8343, 8343, 8343,
  8174, 8332, 7787, 7801, 7811, 7819, 7828, 7833, 7838, 7854, 7854, 7854, 
    7854, 7854, 7854, 8484, 8402, 8402, 8402, 8402, 8402, 8402,
  7685, 7865, 7503, 7520, 7533, 7542, 7553, 7559, 7565, 7585, 7585, 7585, 
    7585, 7585, 7585, 8227, 8263, 8262, 8263, 8263, 8262, 8262,
  7038, 7242, 7209, 7239, 7259, 7275, 7291, 7302, 7312, 7345, 7345, 7345, 
    7345, 7345, 7345, 7969, 8452, 8452, 8452, 8452, 8452, 8452,
  6673, 6897, 6733, 6760, 6779, 6794, 6809, 6819, 6828, 6859, 6859, 6859, 
    6859, 6859, 6859, 7611, 7889, 7889, 7889, 7889, 7889, 7889,
  6109, 6343, 6397, 6426, 6447, 6463, 6478, 6488, 6499, 6532, 6532, 6532, 
    6532, 6532, 6532, 7410, 7735, 7864, 7864, 7864, 7864, 7864,
  5653, 5894, 5775, 5807, 5830, 5848, 5865, 5876, 5889, 5926, 5926, 5926, 
    5926, 5926, 5926, 7086, 7324, 7471, 7471, 7471, 7471, 7471,
  5418, 5708, 5684, 5721, 5748, 5768, 5788, 5801, 5815, 5858, 5858, 5858, 
    5858, 5858, 5858, 7080, 7393, 7546, 7546, 7546, 7546, 7546,
  5497, 5769, 5890, 5925, 5950, 5969, 5987, 5999, 6012, 6053, 6053, 6053, 
    6053, 6053, 6053, 7047, 7477, 7621, 7621, 7621, 7621, 7621,
  5835, 6096, 6155, 6187, 6211, 6228, 6245, 6257, 6269, 6307, 6307, 6307, 
    6307, 6307, 6307, 7291, 7633, 7770, 7770, 7770, 7770, 7770,
  6192, 6436, 6508, 6537, 6558, 6574, 6589, 6599, 6611, 6644, 6644, 6644, 
    6644, 6644, 6644, 7515, 7831, 7957, 7957, 7957, 7957, 7957,
  6542, 6780, 6892, 6919, 6939, 6953, 6967, 6977, 6987, 7018, 7018, 7018, 
    7018, 7018, 7018, 7778, 8086, 8201, 8201, 8201, 8201, 8201,
  6853, 7078, 7110, 7135, 7153, 7166, 7179, 7187, 7197, 7225, 7225, 7225, 
    7225, 7225, 7225, 7994, 8204, 8314, 8314, 8314, 8314, 8314,
  7008, 7204, 7140, 7162, 7177, 7189, 7200, 7208, 7217, 7241, 7241, 7241, 
    7241, 7241, 7241, 8017, 8145, 8252, 8252, 8252, 8252, 8252,
  7136, 7314, 7079, 7099, 7114, 7125, 7135, 7142, 7150, 7173, 7173, 7173, 
    7173, 7173, 7173, 8073, 8061, 8170, 8170, 8170, 8170, 8170,
  7171, 7346, 7141, 7161, 7175, 7185, 7195, 7202, 7210, 7232, 7232, 7232, 
    7232, 7232, 7232, 8082, 8089, 8196, 8196, 8196, 8196, 8196,
  7123, 7310, 7194, 7215, 7230, 7241, 7251, 7258, 7267, 7290, 7290, 7290, 
    7290, 7290, 7290, 8085, 8165, 8271, 8271, 8271, 8271, 8271,
  7067, 7280, 7233, 7256, 7273, 7285, 7297, 7305, 7314, 7340, 7340, 7340, 
    7340, 7340, 7340, 8133, 8257, 8363, 8363, 8363, 8363, 8363,
  6899, 7122, 7081, 7105, 7123, 7136, 7149, 7158, 7168, 7196, 7196, 7196, 
    7196, 7196, 7196, 8038, 8181, 8292, 8292, 8292, 8292, 8292,
  6734, 6957, 6936, 6961, 6979, 6993, 7006, 7015, 7025, 7054, 7054, 7054, 
    7054, 7054, 7054, 7895, 8074, 8188, 8188, 8188, 8188, 8188,
  6456, 6706, 6668, 6697, 6718, 6733, 6749, 6759, 6770, 6803, 6803, 6803, 
    6803, 6803, 6803, 7779, 7965, 8088, 8088, 8088, 8088, 8088,
  6068, 6324, 6220, 6252, 6274, 6291, 6308, 6319, 6331, 6367, 6367, 6367, 
    6367, 6367, 6367, 7488, 7667, 7803, 7803, 7803, 7803, 7803,
  5671, 5944, 5849, 5884, 5908, 5927, 5945, 5958, 5971, 6011, 6011, 6011, 
    6011, 6011, 6011, 7224, 7454, 7601, 7601, 7601, 7601, 7601,
  5282, 5569, 5463, 5501, 5528, 5549, 5569, 5582, 5597, 5640, 5640, 5640, 
    5640, 5640, 5640, 6962, 7224, 7382, 7382, 7382, 7382, 7382,
  5051, 5348, 5269, 5309, 5338, 5359, 5380, 5394, 5409, 5455, 5455, 5455, 
    5455, 5455, 5455, 6808, 7117, 7280, 7280, 7280, 7280, 7280,
  5074, 5374, 5311, 5352, 5380, 5402, 5422, 5437, 5452, 5498, 5498, 5498, 
    5498, 5498, 5498, 6839, 7155, 7318, 7318, 7318, 7318, 7318,
  5404, 5702, 5627, 5666, 5693, 5714, 5734, 5747, 5762, 5806, 5806, 5806, 
    5806, 5806, 5806, 7108, 7373, 7527, 7527, 7527, 7527, 7527,
  6040, 6298, 6328, 6360, 6382, 6399, 6416, 6427, 6439, 6475, 6475, 6475, 
    6475, 6475, 6475, 7458, 7750, 7883, 7883, 7883, 7883, 7883,
  6672, 6887, 7026, 7051, 7068, 7081, 7094, 7102, 7112, 7140, 7140, 7140, 
    7140, 7140, 7140, 7785, 8113, 8223, 8223, 8223, 8223, 8223,
  7235, 7418, 7567, 7586, 7600, 7610, 7620, 7626, 7634, 7655, 7655, 7655, 
    7655, 7655, 7655, 8122, 8404, 8498, 8498, 8498, 8498, 8498,
  7663, 7792, 7835, 7847, 7856, 7862, 7869, 7872, 7878, 7892, 7892, 7892, 
    7892, 7892, 7892, 8268, 8443, 8526, 8526, 8526, 8526, 8526,
  7900, 8038, 8016, 8028, 8037, 8044, 8050, 8054, 8060, 8073, 8073, 8073, 
    8073, 8073, 8073, 8512, 8598, 8677, 8677, 8677, 8677, 8677,
  8010, 8242, 8250, 8253, 8256, 8257, 8259, 8260, 8261, 8264, 8264, 8264, 
    8264, 8264, 8264, 8535, 8381, 8381, 8381, 8381, 8381, 8381,
  7963, 8068, 7996, 8004, 8011, 8016, 8021, 8024, 8028, 8038, 8038, 8038, 
    8038, 8038, 8038, 8435, 8493, 8571, 8571, 8571, 8571, 8571,
  7941, 8067, 8086, 8097, 8105, 8110, 8116, 8119, 8125, 8137, 8137, 8137, 
    8137, 8137, 8137, 8492, 8615, 8692, 8692, 8692, 8692, 8692,
  7999, 8254, 8379, 8373, 8369, 8365, 8362, 8360, 8357, 8350, 8350, 8350, 
    8350, 8350, 8350, 8461, 8113, 8113, 8113, 8113, 8113, 8113,
  8177, 8417, 8533, 8522, 8514, 8508, 8502, 8497, 8493, 8480, 8480, 8480, 
    8480, 8480, 8480, 8495, 8045, 8045, 8045, 8045, 8045, 8045,
  7962, 8214, 8414, 8402, 8393, 8386, 8379, 8374, 8370, 8355, 8355, 8355, 
    8355, 8355, 8355, 8300, 7873, 7873, 7873, 7873, 7873, 7873,
  7700, 7985, 8342, 8326, 8315, 8307, 8299, 8293, 8287, 8269, 8269, 8269, 
    8269, 8269, 8269, 8113, 7680, 7680, 7680, 7680, 7680, 7680,
  7351, 7699, 8199, 8184, 8173, 8165, 8157, 8151, 8146, 8129, 8129, 8129, 
    8129, 8129, 8129, 8018, 7554, 7554, 7554, 7554, 7554, 7555,
  7207, 7617, 8260, 8241, 8229, 8219, 8210, 8203, 8196, 8176, 8176, 8176, 
    8176, 8176, 8176, 8077, 7493, 7493, 7493, 7493, 7493, 7493,
  8617, 8738, 8892, 8895, 8897, 8898, 8901, 8902, 8903, 8906, 8906, 8906, 
    8906, 8906, 8906, 8961, 9031, 9031, 9031, 9031, 9031, 9031,
  8803, 8914, 9069, 9069, 9069, 9069, 9070, 9069, 9069, 9069, 9069, 9069, 
    9069, 9069, 9069, 9068, 9073, 9073, 9073, 9073, 9073, 9073,
  8916, 9025, 9089, 9087, 9085, 9084, 9084, 9083, 9082, 9079, 9079, 9079, 
    9079, 9079, 9079, 9103, 9000, 9000, 9000, 9000, 9000, 9000,
  8921, 9026, 9104, 9099, 9096, 9093, 9091, 9089, 9088, 9082, 9082, 9082, 
    9082, 9082, 9082, 9066, 8905, 8905, 8905, 8905, 8905, 8905,
  9012, 9114, 9064, 9063, 9062, 9061, 9062, 9061, 9061, 9060, 9060, 9060, 
    9060, 9060, 9060, 9125, 9030, 9030, 9030, 9030, 9030, 9030,
  9003, 9102, 9043, 9043, 9043, 9043, 9044, 9044, 9044, 9043, 9043, 9043, 
    9043, 9043, 9043, 9106, 9047, 9047, 9047, 9047, 9047, 9047,
  8980, 9076, 8991, 8988, 8985, 8983, 8982, 8981, 8979, 8975, 8975, 8975, 
    8975, 8975, 8975, 9015, 8850, 8850, 8850, 8850, 8850, 8850,
  9107, 9184, 9104, 9094, 9086, 9081, 9076, 9073, 9069, 9057, 9057, 9057, 
    9057, 9057, 9057, 8973, 8681, 8681, 8681, 8681, 8681, 8681,
  9018, 9113, 8951, 8951, 8950, 8950, 8950, 8950, 8950, 8949, 8949, 8949, 
    8949, 8949, 8949, 9047, 8938, 8938, 8938, 8938, 8938, 8938,
  8975, 9075, 8873, 8875, 8876, 8877, 8879, 8879, 8880, 8881, 8881, 8881, 
    8881, 8881, 8881, 9029, 8952, 8952, 8952, 8952, 8952, 8952,
  8902, 9004, 8888, 8890, 8891, 8892, 8894, 8894, 8895, 8897, 8897, 8897, 
    8897, 8897, 8897, 9011, 8977, 8977, 8977, 8977, 8977, 8977,
  8881, 8985, 8881, 8883, 8885, 8886, 8888, 8889, 8890, 8892, 8892, 8892, 
    8892, 8892, 8892, 9011, 8984, 8984, 8984, 8984, 8984, 8984,
  8923, 9027, 8904, 8905, 8906, 8906, 8908, 8908, 8909, 8910, 8910, 8910, 
    8910, 8910, 8910, 9029, 8966, 8966, 8966, 8966, 8966, 8966,
  8754, 8862, 8643, 8642, 8642, 8641, 8642, 8641, 8641, 8640, 8640, 8640, 
    8640, 8640, 8640, 8811, 8614, 8614, 8614, 8614, 8614, 8614,
  8853, 8963, 8691, 8691, 8690, 8690, 8690, 8690, 8690, 8689, 8689, 8689, 
    8689, 8689, 8689, 8900, 8678, 8678, 8678, 8678, 8678, 8678,
  8657, 8783, 8482, 8486, 8488, 8490, 8493, 8494, 8495, 8499, 8499, 8499, 
    8499, 8499, 8499, 8812, 8638, 8638, 8638, 8638, 8638, 8638,
  8852, 8963, 8643, 8644, 8644, 8645, 8646, 8646, 8647, 8648, 8648, 8648, 
    8648, 8648, 8648, 8899, 8691, 8691, 8691, 8691, 8691, 8691,
  8972, 9072, 8714, 8713, 8713, 8712, 8713, 8713, 8713, 8712, 8712, 8712, 
    8712, 8712, 8712, 8932, 8701, 8701, 8701, 8701, 8701, 8701,
  9005, 9099, 8714, 8712, 8711, 8711, 8711, 8711, 8710, 8709, 8709, 8709, 
    8709, 8709, 8709, 8907, 8670, 8670, 8670, 8670, 8670, 8670,
  8991, 9085, 8826, 8824, 8822, 8821, 8820, 8820, 8819, 8816, 8816, 8816, 
    8816, 8816, 8816, 8942, 8735, 8735, 8735, 8735, 8735, 8735,
  9048, 9142, 8819, 8818, 8817, 8816, 8816, 8816, 8815, 8813, 8813, 8813, 
    8813, 8813, 8813, 8983, 8770, 8770, 8770, 8770, 8770, 8770,
  8975, 9074, 8719, 8719, 8719, 8719, 8720, 8720, 8719, 8719, 8719, 8719, 
    8719, 8719, 8719, 8933, 8721, 8721, 8721, 8721, 8721, 8721,
  8923, 9026, 8626, 8627, 8627, 8627, 8628, 8628, 8629, 8629, 8629, 8629, 
    8629, 8629, 8629, 8886, 8652, 8652, 8652, 8652, 8652, 8652,
  8953, 9058, 8623, 8624, 8625, 8625, 8627, 8627, 8627, 8629, 8629, 8629, 
    8629, 8629, 8629, 8917, 8676, 8676, 8676, 8676, 8676, 8676,
  9015, 9116, 8777, 8776, 8775, 8775, 8775, 8775, 8774, 8773, 8773, 8773, 
    8773, 8773, 8773, 8987, 8750, 8750, 8750, 8750, 8750, 8750,
  9099, 9192, 8834, 8832, 8830, 8828, 8828, 8827, 8826, 8823, 8823, 8823, 
    8823, 8823, 8823, 9001, 8738, 8738, 8738, 8738, 8738, 8738,
  9147, 9236, 8872, 8870, 8869, 8868, 8868, 8867, 8866, 8864, 8864, 8864, 
    8864, 8864, 8864, 9034, 8806, 8806, 8806, 8806, 8806, 8806,
  9253, 9335, 8940, 8938, 8936, 8934, 8934, 8933, 8932, 8929, 8929, 8929, 
    8929, 8929, 8929, 9082, 8843, 8843, 8843, 8843, 8843, 8843,
  9188, 9276, 8877, 8873, 8871, 8869, 8868, 8866, 8865, 8861, 8861, 8861, 
    8861, 8861, 8861, 9033, 8736, 8736, 8736, 8736, 8736, 8736,
  9169, 9269, 8884, 8887, 8890, 8891, 8894, 8895, 8896, 8900, 8900, 8900, 
    8900, 8900, 8900, 9161, 9033, 9033, 9033, 9033, 9033, 9033,
  9060, 9169, 8836, 8841, 8844, 8847, 8850, 8852, 8854, 8859, 8859, 8859, 
    8859, 8859, 8859, 9139, 9053, 9053, 9053, 9053, 9053, 9053,
  8944, 9062, 8689, 8697, 8702, 8706, 8711, 8713, 8716, 8725, 8725, 8725, 
    8725, 8725, 8725, 9078, 9016, 9016, 9016, 9016, 9016, 9016,
  8806, 8933, 8603, 8610, 8616, 8620, 8625, 8627, 8630, 8639, 8639, 8639, 
    8639, 8639, 8639, 9002, 8934, 8934, 8934, 8934, 8934, 8934,
  8744, 8855, 8548, 8549, 8550, 8551, 8553, 8554, 8554, 8556, 8556, 8556, 
    8556, 8556, 8556, 8797, 8624, 8624, 8624, 8624, 8624, 8624,
  8554, 8676, 8403, 8406, 8408, 8410, 8413, 8414, 8415, 8419, 8419, 8419, 
    8419, 8419, 8419, 8697, 8552, 8552, 8552, 8552, 8552, 8552,
  8469, 8597, 8331, 8335, 8338, 8340, 8344, 8345, 8347, 8351, 8351, 8351, 
    8351, 8351, 8351, 8656, 8517, 8517, 8517, 8517, 8517, 8517,
  8373, 8505, 8187, 8192, 8196, 8198, 8202, 8204, 8205, 8211, 8211, 8211, 
    8211, 8211, 8211, 8562, 8405, 8405, 8405, 8405, 8405, 8405,
  8335, 8470, 8226, 8231, 8234, 8237, 8240, 8242, 8244, 8249, 8249, 8249, 
    8249, 8249, 8249, 8576, 8446, 8446, 8446, 8446, 8446, 8446,
  8383, 8508, 8247, 8250, 8252, 8253, 8256, 8257, 8258, 8261, 8261, 8261, 
    8261, 8261, 8261, 8541, 8381, 8381, 8381, 8381, 8381, 8381,
  8305, 8432, 8172, 8173, 8174, 8174, 8176, 8177, 8177, 8178, 8178, 8178, 
    8178, 8178, 8178, 8451, 8234, 8234, 8234, 8234, 8234, 8234,
  8474, 8594, 8264, 8266, 8266, 8267, 8269, 8269, 8270, 8271, 8271, 8271, 
    8271, 8271, 8271, 8557, 8330, 8330, 8330, 8330, 8330, 8330,
  8542, 8659, 8271, 8272, 8272, 8272, 8274, 8274, 8274, 8274, 8274, 8274, 
    8274, 8274, 8274, 8569, 8299, 8299, 8299, 8299, 8299, 8299,
  8471, 8599, 8156, 8156, 8155, 8154, 8155, 8155, 8154, 8153, 8153, 8153, 
    8153, 8153, 8153, 8519, 8130, 8130, 8130, 8130, 8130, 8130,
  8536, 8661, 8376, 8378, 8380, 8382, 8384, 8385, 8386, 8389, 8389, 8389, 
    8389, 8389, 8389, 8685, 8501, 8501, 8501, 8501, 8501, 8501,
  8522, 8648, 8337, 8338, 8339, 8340, 8342, 8342, 8343, 8345, 8345, 8345, 
    8345, 8345, 8345, 8653, 8414, 8414, 8414, 8414, 8414, 8414,
  8606, 8727, 8429, 8430, 8430, 8430, 8431, 8431, 8431, 8432, 8432, 8432, 
    8432, 8432, 8432, 8703, 8452, 8452, 8452, 8452, 8452, 8452,
  8611, 8731, 8569, 8568, 8568, 8567, 8568, 8567, 8567, 8566, 8566, 8566, 
    8566, 8566, 8566, 8756, 8542, 8542, 8542, 8542, 8542, 8542,
  8580, 8703, 8479, 8479, 8478, 8478, 8479, 8479, 8478, 8478, 8478, 8478, 
    8478, 8478, 8478, 8712, 8466, 8466, 8466, 8466, 8466, 8466,
  8700, 8821, 8571, 8572, 8573, 8574, 8576, 8577, 8577, 8579, 8579, 8579, 
    8579, 8579, 8579, 8834, 8643, 8643, 8643, 8643, 8643, 8643,
  8669, 8797, 8486, 8489, 8492, 8494, 8497, 8498, 8500, 8504, 8504, 8504, 
    8504, 8504, 8504, 8836, 8656, 8656, 8656, 8656, 8656, 8656,
  8589, 8710, 8424, 8427, 8429, 8430, 8432, 8433, 8434, 8437, 8437, 8437, 
    8437, 8437, 8437, 8715, 8545, 8545, 8545, 8545, 8545, 8545,
  8593, 8714, 8379, 8382, 8384, 8385, 8388, 8389, 8390, 8393, 8393, 8393, 
    8393, 8393, 8393, 8700, 8511, 8511, 8511, 8511, 8511, 8511,
  8573, 8694, 8435, 8437, 8438, 8438, 8440, 8441, 8441, 8442, 8442, 8442, 
    8442, 8442, 8442, 8698, 8503, 8503, 8503, 8503, 8503, 8503,
  8503, 8629, 8398, 8400, 8402, 8403, 8405, 8406, 8407, 8409, 8409, 8409, 
    8409, 8409, 8409, 8673, 8503, 8503, 8503, 8503, 8503, 8503,
  8532, 8667, 8419, 8421, 8422, 8423, 8425, 8426, 8427, 8429, 8429, 8429, 
    8429, 8429, 8429, 8744, 8511, 8511, 8511, 8511, 8511, 8511,
  8383, 8524, 8150, 8159, 8164, 8169, 8174, 8177, 8180, 8189, 8189, 8189, 
    8189, 8189, 8189, 8630, 8506, 8506, 8506, 8506, 8506, 8506,
  8206, 8353, 7821, 7836, 7847, 7855, 7864, 7870, 7875, 7892, 7892, 7892, 
    7892, 7892, 7892, 8476, 8473, 8473, 8473, 8473, 8473, 8473,
  7934, 8100, 7718, 7732, 7742, 7750, 7758, 7763, 7768, 7784, 7784, 7784, 
    7784, 7784, 7784, 8359, 8327, 8327, 8327, 8327, 8327, 8327,
  7413, 7602, 7484, 7502, 7514, 7523, 7534, 7540, 7546, 7565, 7565, 7565, 
    7565, 7565, 7565, 8108, 8229, 8229, 8229, 8229, 8229, 8229,
  6773, 6993, 6951, 6977, 6995, 7009, 7024, 7033, 7042, 7071, 7071, 7071, 
    7071, 7071, 7071, 7742, 8052, 8052, 8052, 8052, 8052, 8052,
  6457, 6701, 6305, 6338, 6361, 6379, 6397, 6409, 6420, 6457, 6457, 6457, 
    6457, 6457, 6457, 7445, 7697, 7697, 7697, 7697, 7697, 7697,
  5994, 6236, 6176, 6206, 6228, 6245, 6261, 6272, 6284, 6319, 6319, 6319, 
    6319, 6319, 6319, 7370, 7614, 7751, 7751, 7751, 7751, 7751,
  5800, 6062, 6021, 6054, 6078, 6096, 6113, 6125, 6138, 6176, 6176, 6176, 
    6176, 6176, 6176, 7286, 7555, 7698, 7698, 7698, 7698, 7698,
  5803, 6067, 6146, 6179, 6202, 6220, 6237, 6249, 6261, 6299, 6299, 6299, 
    6299, 6299, 6299, 7274, 7635, 7772, 7772, 7772, 7772, 7772,
  6110, 6362, 6414, 6445, 6467, 6483, 6499, 6510, 6522, 6557, 6557, 6557, 
    6557, 6557, 6557, 7486, 7792, 7921, 7921, 7921, 7921, 7921,
  6510, 6742, 6823, 6850, 6869, 6883, 6897, 6906, 6917, 6948, 6948, 6948, 
    6948, 6948, 6948, 7728, 8018, 8135, 8135, 8135, 8135, 8135,
  6772, 6980, 7094, 7117, 7134, 7146, 7159, 7166, 7176, 7202, 7202, 7202, 
    7202, 7202, 7202, 7845, 8140, 8248, 8248, 8248, 8248, 8248,
  7011, 7205, 7235, 7256, 7271, 7283, 7294, 7301, 7310, 7334, 7334, 7334, 
    7334, 7334, 7334, 8000, 8206, 8309, 8309, 8309, 8309, 8309,
  7190, 7373, 7281, 7301, 7315, 7326, 7336, 7343, 7351, 7373, 7373, 7373, 
    7373, 7373, 7373, 8118, 8211, 8314, 8314, 8314, 8314, 8314,
  7296, 7453, 7209, 7226, 7239, 7248, 7257, 7263, 7271, 7291, 7291, 7291, 
    7291, 7291, 7291, 8125, 8099, 8204, 8204, 8204, 8204, 8204,
  7306, 7471, 7317, 7335, 7348, 7357, 7367, 7373, 7380, 7400, 7400, 7400, 
    7400, 7400, 7400, 8148, 8186, 8288, 8288, 8288, 8288, 8288,
  7302, 7479, 7440, 7458, 7472, 7482, 7492, 7498, 7505, 7527, 7527, 7527, 
    7527, 7527, 7527, 8179, 8304, 8402, 8402, 8402, 8402, 8402,
  7249, 7441, 7383, 7404, 7418, 7429, 7440, 7447, 7455, 7478, 7478, 7478, 
    7478, 7478, 7478, 8203, 8307, 8407, 8407, 8407, 8407, 8407,
  7122, 7325, 7255, 7277, 7293, 7304, 7316, 7323, 7332, 7357, 7357, 7357, 
    7357, 7357, 7357, 8142, 8244, 8348, 8348, 8348, 8348, 8348,
  6893, 7117, 7063, 7088, 7106, 7120, 7133, 7141, 7151, 7179, 7179, 7179, 
    7179, 7179, 7179, 8040, 8174, 8286, 8286, 8286, 8286, 8286,
  6691, 6933, 6933, 6960, 6980, 6994, 7009, 7018, 7029, 7060, 7060, 7060, 
    7060, 7060, 7060, 7938, 8131, 8247, 8247, 8247, 8247, 8247,
  6360, 6622, 6579, 6610, 6632, 6648, 6665, 6675, 6687, 6722, 6722, 6722, 
    6722, 6722, 6722, 7753, 7941, 8068, 8068, 8068, 8068, 8068,
  5934, 6208, 6095, 6129, 6154, 6172, 6190, 6201, 6215, 6254, 6254, 6254, 
    6254, 6254, 6254, 7454, 7635, 7776, 7776, 7776, 7776, 7776,
  5518, 5808, 5638, 5676, 5703, 5723, 5742, 5755, 5770, 5813, 5813, 5813, 
    5813, 5813, 5813, 7180, 7358, 7512, 7512, 7512, 7512, 7512,
  5273, 5576, 5420, 5460, 5488, 5510, 5531, 5545, 5560, 5606, 5606, 5606, 
    5606, 5606, 5606, 7032, 7244, 7405, 7405, 7405, 7405, 7405,
  5292, 5589, 5426, 5465, 5493, 5514, 5534, 5548, 5563, 5608, 5608, 5608, 
    5608, 5608, 5608, 7021, 7228, 7388, 7388, 7388, 7388, 7388,
  5651, 5928, 5769, 5804, 5830, 5849, 5867, 5880, 5894, 5935, 5935, 5935, 
    5935, 5935, 5935, 7236, 7412, 7562, 7562, 7562, 7562, 7562,
  6185, 6428, 6388, 6418, 6439, 6455, 6471, 6481, 6493, 6527, 6527, 6527, 
    6527, 6527, 6527, 7523, 7749, 7879, 7879, 7879, 7879, 7879,
  6706, 6910, 6962, 6986, 7003, 7015, 7028, 7036, 7045, 7072, 7072, 7072, 
    7072, 7072, 7072, 7782, 8041, 8152, 8152, 8152, 8152, 8152,
  7309, 7484, 7566, 7583, 7597, 7606, 7616, 7621, 7629, 7649, 7649, 7649, 
    7649, 7649, 7649, 8157, 8380, 8473, 8473, 8473, 8473, 8473,
  7785, 7949, 8001, 8016, 8027, 8035, 8043, 8047, 8054, 8071, 8071, 8071, 
    8071, 8071, 8071, 8515, 8660, 8742, 8742, 8742, 8742, 8742,
  7908, 8033, 8003, 8013, 8022, 8028, 8034, 8037, 8042, 8054, 8054, 8054, 
    8054, 8054, 8054, 8468, 8553, 8633, 8633, 8633, 8633, 8633,
  7945, 8059, 7945, 7955, 7962, 7968, 7973, 7976, 7981, 7993, 7993, 7993, 
    7993, 7993, 7993, 8465, 8488, 8569, 8569, 8569, 8569, 8569,
  8038, 8230, 8220, 8222, 8223, 8224, 8225, 8225, 8226, 8228, 8228, 8228, 
    8228, 8228, 8228, 8373, 8288, 8288, 8288, 8288, 8288, 8288,
  8057, 8197, 8242, 8253, 8262, 8268, 8274, 8278, 8283, 8296, 8296, 8296, 
    8296, 8296, 8296, 8642, 8764, 8838, 8838, 8838, 8838, 8838,
  8137, 8337, 8346, 8342, 8339, 8337, 8335, 8333, 8331, 8327, 8327, 8327, 
    8327, 8327, 8327, 8418, 8174, 8174, 8174, 8174, 8174, 8174,
  8199, 8383, 8403, 8394, 8388, 8383, 8378, 8375, 8371, 8362, 8362, 8362, 
    8362, 8362, 8362, 8331, 8022, 8022, 8022, 8022, 8022, 8022,
  7996, 8202, 8327, 8316, 8308, 8302, 8296, 8292, 8287, 8275, 8275, 8275, 
    8275, 8275, 8275, 8176, 7850, 7850, 7850, 7850, 7850, 7850,
  7854, 8135, 8467, 8449, 8437, 8427, 8417, 8411, 8404, 8384, 8384, 8384, 
    8384, 8384, 8384, 8217, 7700, 7700, 7700, 7700, 7700, 7700,
  7601, 7943, 8421, 8404, 8392, 8384, 8375, 8368, 8362, 8344, 8344, 8344, 
    8344, 8344, 8344, 8226, 7714, 7714, 7714, 7714, 7714, 7714,
  7395, 7757, 8300, 8284, 8274, 8266, 8257, 8252, 8246, 8228, 8228, 8228, 
    8228, 8228, 8228, 8112, 7643, 7643, 7643, 7643, 7643, 7644,
  8627, 8746, 8947, 8950, 8951, 8953, 8955, 8955, 8956, 8959, 8959, 8959, 
    8959, 8959, 8959, 8980, 9058, 9058, 9058, 9058, 9058, 9058,
  8855, 8964, 8965, 8965, 8965, 8965, 8966, 8966, 8966, 8966, 8966, 8966, 
    8966, 8966, 8966, 9041, 8979, 8979, 8979, 8979, 8979, 8979,
  8918, 9022, 8989, 8988, 8987, 8987, 8987, 8987, 8986, 8985, 8985, 8985, 
    8985, 8985, 8985, 9049, 8956, 8956, 8955, 8955, 8956, 8956,
  9029, 9128, 9103, 9100, 9097, 9095, 9094, 9092, 9091, 9087, 9087, 9087, 
    9087, 9087, 9087, 9110, 8953, 8953, 8953, 8953, 8953, 8953,
  9005, 9103, 9175, 9170, 9167, 9164, 9162, 9161, 9159, 9153, 9153, 9153, 
    9153, 9153, 9153, 9117, 8983, 8983, 8983, 8983, 8983, 8983,
  9002, 9099, 9050, 9047, 9045, 9043, 9042, 9041, 9040, 9036, 9036, 9036, 
    9036, 9036, 9036, 9066, 8923, 8923, 8923, 8923, 8923, 8923,
  9107, 9187, 9149, 9140, 9133, 9128, 9124, 9121, 9118, 9107, 9107, 9107, 
    9107, 9107, 9107, 9023, 8766, 8766, 8766, 8766, 8766, 8766,
  9005, 9091, 8940, 8936, 8933, 8930, 8929, 8927, 8926, 8921, 8921, 8921, 
    8921, 8921, 8921, 8945, 8769, 8769, 8769, 8769, 8769, 8769,
  8970, 9069, 8933, 8934, 8934, 8934, 8935, 8935, 8936, 8936, 8936, 8936, 
    8936, 8936, 8936, 9038, 8959, 8959, 8959, 8959, 8959, 8959,
  9006, 9104, 8927, 8928, 8929, 8929, 8931, 8931, 8932, 8933, 8933, 8933, 
    8933, 8933, 8933, 9060, 8987, 8987, 8987, 8987, 8987, 8987,
  8933, 9033, 8909, 8910, 8910, 8911, 8912, 8913, 8913, 8914, 8914, 8914, 
    8914, 8914, 8914, 9016, 8963, 8963, 8963, 8963, 8963, 8963,
  8862, 8966, 8846, 8846, 8847, 8847, 8848, 8848, 8849, 8849, 8849, 8849, 
    8849, 8849, 8849, 8964, 8881, 8881, 8881, 8881, 8881, 8881,
  8792, 8893, 8651, 8648, 8646, 8644, 8644, 8643, 8642, 8638, 8638, 8638, 
    8638, 8638, 8638, 8776, 8532, 8532, 8532, 8532, 8532, 8532,
  9035, 9121, 8921, 8911, 8905, 8900, 8896, 8892, 8889, 8878, 8878, 8878, 
    8878, 8878, 8878, 8899, 8530, 8530, 8530, 8530, 8530, 8530,
  8878, 8984, 8721, 8720, 8720, 8719, 8720, 8720, 8719, 8718, 8718, 8718, 
    8718, 8718, 8718, 8907, 8699, 8699, 8699, 8699, 8699, 8699,
  8926, 9030, 8714, 8714, 8713, 8713, 8714, 8714, 8714, 8713, 8713, 8713, 
    8713, 8713, 8713, 8924, 8705, 8705, 8705, 8705, 8705, 8705,
  9053, 9139, 8833, 8827, 8823, 8819, 8817, 8815, 8813, 8807, 8807, 8807, 
    8807, 8807, 8807, 8910, 8599, 8599, 8599, 8599, 8599, 8599,
  8824, 8936, 8540, 8542, 8543, 8543, 8545, 8545, 8546, 8547, 8547, 8547, 
    8547, 8547, 8547, 8840, 8607, 8607, 8607, 8607, 8607, 8607,
  8852, 8958, 8652, 8652, 8652, 8653, 8654, 8654, 8654, 8654, 8654, 8654, 
    8654, 8654, 8654, 8868, 8671, 8671, 8671, 8671, 8671, 8671,
  8964, 9065, 8689, 8689, 8689, 8689, 8690, 8690, 8690, 8690, 8690, 8690, 
    8690, 8690, 8690, 8922, 8696, 8696, 8696, 8696, 8696, 8696,
  8921, 9023, 8653, 8653, 8653, 8653, 8654, 8654, 8654, 8654, 8654, 8654, 
    8654, 8654, 8654, 8889, 8666, 8666, 8666, 8666, 8666, 8666,
  8995, 9092, 8735, 8735, 8734, 8734, 8735, 8735, 8735, 8734, 8734, 8734, 
    8734, 8734, 8734, 8938, 8734, 8734, 8734, 8734, 8734, 8734,
  9012, 9109, 8713, 8713, 8713, 8713, 8713, 8713, 8713, 8713, 8713, 8713, 
    8713, 8713, 8713, 8937, 8711, 8711, 8711, 8711, 8711, 8711,
  8931, 9036, 8604, 8604, 8603, 8603, 8604, 8604, 8603, 8603, 8603, 8603, 
    8603, 8603, 8603, 8874, 8597, 8597, 8597, 8597, 8597, 8597,
  8908, 9017, 8572, 8573, 8574, 8575, 8576, 8577, 8577, 8578, 8578, 8578, 
    8578, 8578, 8578, 8885, 8631, 8631, 8631, 8631, 8631, 8631,
  8941, 9047, 8617, 8618, 8618, 8618, 8620, 8620, 8620, 8621, 8621, 8621, 
    8621, 8621, 8621, 8904, 8650, 8650, 8650, 8650, 8650, 8650,
  9110, 9205, 9022, 9019, 9017, 9015, 9015, 9014, 9013, 9010, 9010, 9010, 
    9010, 9010, 9010, 9104, 8913, 8913, 8913, 8913, 8913, 8913,
  9188, 9272, 8893, 8891, 8889, 8888, 8888, 8888, 8887, 8885, 8885, 8885, 
    8885, 8885, 8885, 9043, 8822, 8822, 8822, 8822, 8822, 8822,
  9240, 9336, 9041, 9043, 9044, 9044, 9046, 9047, 9047, 9049, 9049, 9049, 
    9049, 9049, 9049, 9237, 9119, 9119, 9119, 9119, 9119, 9119,
  9108, 9215, 8968, 8969, 8969, 8970, 8971, 8972, 8972, 8973, 8973, 8973, 
    8973, 8973, 8973, 9175, 9019, 9019, 9019, 9019, 9019, 9019,
  8994, 9107, 8813, 8814, 8814, 8815, 8816, 8817, 8817, 8818, 8818, 8818, 
    8818, 8818, 8818, 9069, 8865, 8865, 8865, 8865, 8865, 8865,
  8955, 9072, 8838, 8842, 8845, 8847, 8850, 8851, 8853, 8857, 8857, 8857, 
    8857, 8857, 8857, 9110, 9011, 9011, 9011, 9011, 9011, 9011,
  8808, 8934, 8597, 8605, 8611, 8615, 8621, 8623, 8626, 8636, 8636, 8636, 
    8636, 8636, 8636, 9005, 8956, 8956, 8956, 8956, 8956, 8956,
  8811, 8918, 8567, 8568, 8569, 8569, 8571, 8571, 8571, 8572, 8572, 8572, 
    8572, 8572, 8572, 8820, 8616, 8616, 8616, 8616, 8616, 8616,
  8726, 8837, 8552, 8553, 8553, 8553, 8555, 8555, 8555, 8556, 8556, 8556, 
    8556, 8556, 8556, 8780, 8591, 8591, 8591, 8591, 8591, 8591,
  8681, 8797, 8448, 8450, 8452, 8454, 8456, 8457, 8458, 8461, 8461, 8461, 
    8461, 8461, 8461, 8755, 8571, 8571, 8571, 8571, 8571, 8571,
  8627, 8744, 8400, 8403, 8405, 8406, 8409, 8410, 8411, 8414, 8414, 8414, 
    8414, 8414, 8414, 8712, 8537, 8537, 8537, 8537, 8537, 8537,
  8586, 8709, 8211, 8214, 8217, 8219, 8222, 8223, 8224, 8228, 8228, 8228, 
    8228, 8228, 8228, 8633, 8374, 8374, 8374, 8374, 8374, 8374,
  8605, 8721, 8283, 8286, 8287, 8288, 8291, 8292, 8292, 8295, 8295, 8295, 
    8295, 8295, 8295, 8631, 8394, 8394, 8394, 8394, 8394, 8394,
  8654, 8765, 8492, 8493, 8494, 8494, 8496, 8496, 8496, 8497, 8497, 8497, 
    8497, 8497, 8497, 8717, 8536, 8536, 8536, 8536, 8536, 8536,
  8420, 8543, 8173, 8177, 8180, 8182, 8185, 8187, 8188, 8192, 8192, 8192, 
    8192, 8192, 8192, 8529, 8351, 8351, 8351, 8351, 8351, 8351,
  8555, 8680, 8324, 8324, 8324, 8324, 8325, 8325, 8325, 8325, 8325, 8325, 
    8325, 8325, 8325, 8639, 8332, 8332, 8332, 8332, 8332, 8332,
  8549, 8675, 8271, 8272, 8273, 8274, 8276, 8276, 8277, 8278, 8278, 8278, 
    8278, 8278, 8278, 8632, 8346, 8346, 8346, 8346, 8346, 8346,
  8616, 8742, 8364, 8365, 8366, 8366, 8367, 8368, 8368, 8369, 8369, 8369, 
    8369, 8369, 8369, 8705, 8407, 8407, 8407, 8407, 8407, 8407,
  8693, 8811, 8497, 8497, 8497, 8497, 8499, 8499, 8499, 8499, 8499, 8499, 
    8499, 8499, 8499, 8770, 8519, 8519, 8519, 8519, 8519, 8519,
  8760, 8871, 8598, 8594, 8591, 8589, 8588, 8587, 8585, 8581, 8581, 8581, 
    8581, 8581, 8581, 8775, 8449, 8449, 8449, 8449, 8449, 8449,
  8828, 8935, 8768, 8762, 8758, 8755, 8753, 8751, 8748, 8741, 8741, 8741, 
    8741, 8741, 8741, 8854, 8525, 8525, 8525, 8525, 8525, 8525,
  8833, 8940, 8753, 8746, 8741, 8737, 8735, 8732, 8730, 8722, 8722, 8722, 
    8722, 8722, 8722, 8840, 8476, 8476, 8476, 8476, 8476, 8476,
  8788, 8903, 8707, 8704, 8703, 8701, 8701, 8700, 8699, 8696, 8696, 8696, 
    8696, 8696, 8696, 8881, 8604, 8604, 8604, 8604, 8604, 8604,
  8774, 8893, 8673, 8673, 8674, 8674, 8675, 8675, 8676, 8676, 8676, 8676, 
    8676, 8676, 8676, 8905, 8708, 8708, 8708, 8708, 8708, 8708,
  8825, 8943, 8679, 8680, 8681, 8681, 8683, 8683, 8684, 8685, 8685, 8685, 
    8685, 8685, 8685, 8937, 8732, 8732, 8732, 8732, 8732, 8732,
  8848, 8966, 8712, 8711, 8711, 8711, 8711, 8711, 8711, 8710, 8710, 8710, 
    8710, 8710, 8710, 8951, 8701, 8701, 8701, 8701, 8701, 8701,
  8782, 8895, 8701, 8698, 8696, 8694, 8693, 8692, 8691, 8687, 8687, 8687, 
    8687, 8687, 8687, 8857, 8574, 8574, 8574, 8574, 8574, 8574,
  8632, 8750, 8637, 8639, 8641, 8642, 8644, 8645, 8646, 8648, 8648, 8648, 
    8648, 8648, 8648, 8827, 8743, 8743, 8743, 8743, 8743, 8743,
  8554, 8679, 8459, 8463, 8466, 8468, 8472, 8473, 8475, 8480, 8480, 8480, 
    8480, 8480, 8480, 8753, 8651, 8651, 8651, 8651, 8651, 8651,
  8497, 8623, 8424, 8425, 8426, 8427, 8428, 8429, 8429, 8431, 8431, 8431, 
    8431, 8431, 8431, 8679, 8495, 8495, 8495, 8495, 8495, 8495,
  8238, 8385, 8052, 8069, 8081, 8090, 8100, 8106, 8112, 8131, 8131, 8131, 
    8131, 8131, 8131, 8629, 8782, 8782, 8782, 8782, 8782, 8782,
  7946, 8112, 7705, 7730, 7748, 7761, 7775, 7784, 7793, 7821, 7821, 7821, 
    7821, 7821, 7821, 8478, 8769, 8769, 8769, 8769, 8769, 8769,
  7620, 7796, 7509, 7529, 7543, 7554, 7565, 7572, 7579, 7602, 7602, 7602, 
    7602, 7602, 7602, 8197, 8364, 8364, 8364, 8364, 8364, 8364,
  7029, 7241, 7129, 7150, 7166, 7177, 7190, 7197, 7205, 7229, 7229, 7229, 
    7229, 7229, 7229, 7882, 8052, 8052, 8052, 8052, 8052, 8052,
  6605, 6841, 6485, 6515, 6537, 6553, 6570, 6581, 6592, 6626, 6626, 6626, 
    6626, 6626, 6626, 7551, 7779, 7779, 7779, 7779, 7779, 7779,
  6295, 6529, 6453, 6481, 6502, 6517, 6532, 6542, 6553, 6586, 6586, 6586, 
    6586, 6586, 6586, 7585, 7779, 7908, 7908, 7908, 7908, 7908,
  6095, 6339, 6296, 6327, 6348, 6365, 6380, 6391, 6403, 6438, 6438, 6438, 
    6438, 6438, 6438, 7455, 7697, 7831, 7831, 7831, 7831, 7831,
  6184, 6450, 6518, 6549, 6572, 6589, 6605, 6616, 6628, 6664, 6664, 6664, 
    6664, 6664, 6664, 7603, 7904, 8033, 8033, 8033, 8033, 8033,
  6463, 6698, 6747, 6774, 6794, 6809, 6823, 6833, 6844, 6875, 6875, 6875, 
    6875, 6875, 6875, 7713, 7980, 8099, 8099, 8099, 8099, 8099,
  6788, 7018, 7103, 7128, 7146, 7160, 7173, 7182, 7192, 7221, 7221, 7221, 
    7221, 7221, 7221, 7955, 8212, 8322, 8322, 8322, 8322, 8322,
  6978, 7178, 7286, 7307, 7323, 7335, 7346, 7353, 7362, 7386, 7386, 7386, 
    7386, 7386, 7386, 7981, 8252, 8354, 8354, 8354, 8354, 8354,
  7214, 7414, 7448, 7468, 7484, 7495, 7506, 7513, 7522, 7545, 7545, 7545, 
    7545, 7545, 7545, 8195, 8377, 8476, 8476, 8476, 8476, 8476,
  7354, 7530, 7455, 7473, 7487, 7497, 7506, 7512, 7520, 7541, 7541, 7541, 
    7541, 7541, 7541, 8224, 8314, 8413, 8413, 8413, 8413, 8413,
  7426, 7589, 7421, 7438, 7451, 7460, 7469, 7475, 7482, 7502, 7502, 7502, 
    7502, 7502, 7502, 8247, 8263, 8363, 8363, 8363, 8363, 8363,
  7438, 7607, 7598, 7615, 7627, 7636, 7646, 7651, 7658, 7678, 7678, 7678, 
    7678, 7678, 7678, 8258, 8393, 8485, 8485, 8485, 8485, 8485,
  7404, 7585, 7582, 7600, 7613, 7623, 7633, 7639, 7646, 7667, 7667, 7667, 
    7667, 7667, 7667, 8274, 8409, 8503, 8503, 8503, 8503, 8503,
  7337, 7531, 7499, 7519, 7533, 7544, 7555, 7561, 7570, 7592, 7592, 7592, 
    7592, 7592, 7592, 8282, 8395, 8493, 8493, 8493, 8493, 8493,
  7210, 7411, 7351, 7372, 7387, 7399, 7410, 7417, 7426, 7450, 7450, 7450, 
    7450, 7450, 7450, 8207, 8309, 8412, 8412, 8412, 8412, 8412,
  7071, 7290, 7267, 7290, 7307, 7320, 7332, 7340, 7349, 7376, 7376, 7376, 
    7376, 7376, 7376, 8161, 8301, 8407, 8407, 8407, 8407, 8407,
  6912, 7143, 7133, 7158, 7177, 7190, 7203, 7212, 7222, 7251, 7251, 7251, 
    7251, 7251, 7251, 8075, 8237, 8347, 8347, 8347, 8347, 8347,
  6602, 6850, 6868, 6896, 6916, 6932, 6946, 6956, 6967, 6999, 6999, 6999, 
    6999, 6999, 6999, 7887, 8102, 8220, 8220, 8220, 8220, 8220,
  6242, 6497, 6374, 6405, 6427, 6444, 6460, 6470, 6482, 6518, 6518, 6518, 
    6518, 6518, 6518, 7632, 7775, 7907, 7907, 7907, 7907, 7907,
  5894, 6149, 5884, 5917, 5941, 5958, 5975, 5987, 6000, 6038, 6038, 6038, 
    6038, 6038, 6038, 7362, 7437, 7583, 7583, 7583, 7583, 7583,
  5643, 5902, 5578, 5612, 5637, 5656, 5673, 5686, 5699, 5739, 5739, 5739, 
    5739, 5739, 5739, 7177, 7234, 7389, 7389, 7389, 7389, 7389,
  5620, 5874, 5590, 5624, 5648, 5667, 5684, 5696, 5709, 5749, 5749, 5749, 
    5749, 5749, 5749, 7134, 7229, 7383, 7383, 7383, 7383, 7383,
  5887, 6119, 5994, 6025, 6046, 6063, 6078, 6089, 6101, 6136, 6136, 6136, 
    6136, 6136, 6136, 7239, 7444, 7585, 7585, 7585, 7585, 7585,
  6315, 6513, 6402, 6427, 6445, 6459, 6472, 6480, 6491, 6520, 6520, 6520, 
    6520, 6520, 6520, 7451, 7636, 7763, 7763, 7763, 7763, 7763,
  6899, 7090, 7077, 7098, 7114, 7125, 7137, 7144, 7153, 7178, 7178, 7178, 
    7178, 7178, 7178, 7900, 8089, 8197, 8197, 8197, 8197, 8197,
  7326, 7479, 7550, 7566, 7577, 7586, 7594, 7599, 7606, 7624, 7624, 7624, 
    7624, 7624, 7624, 8082, 8308, 8400, 8400, 8400, 8400, 8400,
  7731, 7880, 7894, 7907, 7918, 7925, 7932, 7937, 7943, 7959, 7959, 7959, 
    7959, 7959, 7959, 8411, 8542, 8626, 8626, 8626, 8626, 8626,
  7898, 8027, 7927, 7939, 7947, 7954, 7960, 7963, 7969, 7982, 7982, 7982, 
    7982, 7982, 7982, 8485, 8512, 8594, 8594, 8594, 8594, 8594,
  7972, 8090, 8109, 8118, 8126, 8131, 8137, 8139, 8144, 8155, 8155, 8155, 
    8155, 8155, 8155, 8484, 8608, 8683, 8683, 8683, 8683, 8683,
  8003, 8131, 8112, 8122, 8130, 8136, 8142, 8145, 8150, 8162, 8162, 8162, 
    8162, 8162, 8162, 8555, 8637, 8714, 8714, 8714, 8714, 8714,
  8041, 8144, 8109, 8117, 8124, 8128, 8132, 8135, 8139, 8149, 8149, 8149, 
    8149, 8149, 8149, 8486, 8567, 8643, 8643, 8643, 8643, 8643,
  8096, 8287, 8291, 8286, 8282, 8279, 8277, 8274, 8272, 8267, 8267, 8267, 
    8267, 8267, 8267, 8316, 8066, 8066, 8066, 8066, 8066, 8066,
  8174, 8369, 8455, 8443, 8435, 8428, 8422, 8417, 8413, 8399, 8399, 8399, 
    8399, 8399, 8399, 8294, 7942, 7942, 7942, 7942, 7942, 7942,
  8140, 8362, 8497, 8483, 8474, 8467, 8460, 8455, 8450, 8435, 8435, 8435, 
    8435, 8435, 8435, 8352, 7930, 7930, 7930, 7930, 7930, 7930,
  7967, 8245, 8543, 8525, 8513, 8503, 8494, 8487, 8480, 8460, 8460, 8460, 
    8460, 8460, 8460, 8324, 7782, 7782, 7782, 7782, 7782, 7782,
  7763, 8105, 8563, 8542, 8528, 8517, 8506, 8498, 8490, 8467, 8467, 8467, 
    8467, 8467, 8467, 8325, 7682, 7682, 7682, 7682, 7682, 7682,
  7621, 7994, 8547, 8524, 8508, 8496, 8484, 8476, 8468, 8442, 8442, 8442, 
    8442, 8442, 8442, 8276, 7590, 7589, 7589, 7589, 7590, 7590,
  8646, 8767, 9022, 9022, 9022, 9022, 9023, 9023, 9023, 9023, 9023, 9023, 
    9023, 9023, 9023, 9007, 9028, 9028, 9028, 9028, 9028, 9028,
  8731, 8845, 9032, 9031, 9029, 9028, 9029, 9028, 9027, 9025, 9025, 9025, 
    9025, 9025, 9025, 9006, 8973, 8973, 8973, 8973, 8973, 8973,
  8885, 8989, 9125, 9121, 9119, 9117, 9116, 9115, 9114, 9110, 9110, 9110, 
    9110, 9110, 9110, 9067, 8991, 8991, 8991, 8991, 8991, 8991,
  8970, 9069, 9063, 9060, 9057, 9056, 9055, 9053, 9052, 9048, 9048, 9048, 
    9048, 9048, 9048, 9066, 8930, 8930, 8930, 8930, 8930, 8930,
  8989, 9085, 9041, 9038, 9036, 9035, 9034, 9033, 9032, 9029, 9029, 9029, 
    9029, 9029, 9029, 9057, 8935, 8935, 8935, 8935, 8935, 8935,
  9184, 9273, 9284, 9269, 9259, 9251, 9244, 9239, 9234, 9217, 9217, 9217, 
    9217, 9217, 9217, 9119, 8674, 8674, 8674, 8674, 8674, 8674,
  9192, 9263, 9217, 9205, 9197, 9191, 9186, 9181, 9177, 9164, 9164, 9164, 
    9164, 9164, 9164, 9033, 8732, 8732, 8732, 8732, 8732, 8732,
  9150, 9221, 9046, 9037, 9031, 9026, 9023, 9020, 9017, 9007, 9007, 9007, 
    9007, 9007, 9007, 8955, 8689, 8689, 8689, 8689, 8689, 8689,
  8971, 9071, 8953, 8954, 8955, 8955, 8956, 8957, 8957, 8958, 8958, 8958, 
    8958, 8958, 8958, 9057, 9000, 9000, 9000, 9000, 9000, 9000,
  8958, 9058, 8923, 8924, 8925, 8925, 8927, 8927, 8927, 8928, 8928, 8928, 
    8928, 8928, 8928, 9040, 8978, 8978, 8978, 8978, 8978, 8978,
  8888, 8992, 8887, 8889, 8890, 8890, 8892, 8892, 8893, 8894, 8894, 8894, 
    8894, 8894, 8894, 9009, 8953, 8953, 8953, 8953, 8953, 8953,
  8893, 8998, 8926, 8927, 8927, 8927, 8929, 8929, 8929, 8930, 8930, 8930, 
    8930, 8930, 8930, 9028, 8970, 8970, 8970, 8970, 8970, 8970,
  8629, 8741, 8544, 8543, 8543, 8542, 8543, 8543, 8543, 8542, 8542, 8542, 
    8542, 8542, 8542, 8717, 8529, 8529, 8529, 8529, 8529, 8529,
  9009, 9100, 8928, 8918, 8911, 8905, 8901, 8898, 8894, 8882, 8882, 8882, 
    8882, 8882, 8882, 8905, 8511, 8511, 8511, 8511, 8511, 8511,
  9002, 9095, 8864, 8861, 8858, 8856, 8855, 8854, 8853, 8849, 8849, 8849, 
    8849, 8849, 8849, 8957, 8730, 8730, 8730, 8730, 8730, 8730,
  9123, 9208, 8957, 8951, 8947, 8944, 8942, 8940, 8938, 8931, 8931, 8931, 
    8931, 8931, 8931, 8998, 8719, 8719, 8719, 8719, 8719, 8719,
  8787, 8901, 8606, 8607, 8608, 8609, 8611, 8611, 8611, 8613, 8613, 8613, 
    8613, 8613, 8613, 8867, 8673, 8673, 8673, 8673, 8673, 8673,
  8885, 8993, 8652, 8653, 8653, 8654, 8655, 8655, 8656, 8657, 8657, 8657, 
    8657, 8657, 8657, 8903, 8696, 8696, 8696, 8696, 8696, 8696,
  8941, 9041, 8711, 8711, 8710, 8710, 8710, 8710, 8710, 8709, 8709, 8709, 
    8709, 8709, 8709, 8910, 8695, 8695, 8695, 8695, 8695, 8695,
  9048, 9144, 8820, 8817, 8814, 8813, 8812, 8811, 8810, 8807, 8807, 8807, 
    8807, 8807, 8807, 8973, 8704, 8704, 8704, 8704, 8704, 8704,
  8946, 9047, 8708, 8708, 8707, 8707, 8708, 8708, 8708, 8707, 8707, 8707, 
    8707, 8707, 8707, 8918, 8706, 8706, 8706, 8706, 8706, 8706,
  9079, 9169, 8789, 8788, 8788, 8787, 8788, 8787, 8787, 8786, 8786, 8786, 
    8786, 8786, 8786, 8972, 8765, 8765, 8765, 8765, 8765, 8765,
  8429, 8553, 8220, 8224, 8226, 8228, 8231, 8233, 8234, 8238, 8238, 8238, 
    8238, 8238, 8238, 8556, 8389, 8389, 8389, 8389, 8389, 8389,
  8840, 8945, 8463, 8464, 8464, 8465, 8466, 8466, 8467, 8467, 8467, 8467, 
    8467, 8467, 8467, 8772, 8505, 8505, 8505, 8505, 8505, 8505,
  8777, 8888, 8509, 8511, 8512, 8513, 8514, 8515, 8515, 8517, 8517, 8517, 
    8517, 8517, 8517, 8797, 8581, 8581, 8581, 8581, 8581, 8581,
  8906, 9007, 8688, 8687, 8686, 8686, 8686, 8686, 8685, 8684, 8684, 8684, 
    8684, 8684, 8684, 8883, 8657, 8657, 8657, 8657, 8657, 8657,
  9044, 9136, 8791, 8790, 8789, 8788, 8789, 8788, 8788, 8787, 8787, 8787, 
    8787, 8787, 8787, 8960, 8754, 8754, 8754, 8754, 8754, 8754,
  9044, 9134, 8751, 8749, 8748, 8748, 8748, 8747, 8747, 8745, 8745, 8745, 
    8745, 8745, 8745, 8931, 8702, 8702, 8702, 8702, 8702, 8702,
  9092, 9193, 8898, 8900, 8901, 8902, 8903, 8904, 8904, 8906, 8906, 8906, 
    8906, 8906, 8906, 9113, 8970, 8970, 8970, 8970, 8970, 8970,
  8954, 9063, 8763, 8766, 8768, 8769, 8772, 8773, 8774, 8777, 8777, 8777, 
    8777, 8777, 8777, 9020, 8887, 8887, 8887, 8887, 8887, 8887,
  9024, 9138, 8766, 8774, 8779, 8783, 8789, 8791, 8794, 8803, 8803, 8803, 
    8803, 8803, 8803, 9140, 9108, 9108, 9108, 9108, 9108, 9108,
  8915, 9030, 8640, 8648, 8653, 8657, 8663, 8665, 8668, 8677, 8677, 8677, 
    8677, 8677, 8677, 9028, 8981, 8981, 8981, 8981, 8981, 8981,
  8893, 9009, 8658, 8664, 8668, 8671, 8675, 8677, 8679, 8685, 8685, 8685, 
    8685, 8685, 8685, 9001, 8901, 8901, 8901, 8901, 8901, 8901,
  8914, 9014, 8694, 8692, 8690, 8689, 8689, 8688, 8687, 8685, 8685, 8685, 
    8685, 8685, 8685, 8867, 8611, 8611, 8611, 8611, 8611, 8611,
  8800, 8921, 8525, 8532, 8537, 8541, 8546, 8548, 8551, 8559, 8559, 8559, 
    8559, 8559, 8559, 8928, 8836, 8836, 8836, 8836, 8836, 8836,
  8716, 8832, 8404, 8406, 8408, 8410, 8412, 8413, 8414, 8417, 8417, 8417, 
    8417, 8417, 8417, 8747, 8528, 8528, 8528, 8528, 8528, 8528,
  8664, 8789, 8351, 8357, 8361, 8364, 8369, 8371, 8373, 8379, 8379, 8379, 
    8379, 8379, 8379, 8776, 8611, 8611, 8611, 8611, 8611, 8611,
  8729, 8848, 8358, 8363, 8366, 8368, 8372, 8373, 8375, 8380, 8380, 8380, 
    8380, 8380, 8380, 8771, 8558, 8558, 8558, 8558, 8558, 8558,
  8739, 8842, 8332, 8332, 8332, 8332, 8333, 8333, 8333, 8333, 8333, 8333, 
    8333, 8333, 8333, 8637, 8342, 8342, 8342, 8342, 8342, 8342,
  8729, 8834, 8434, 8433, 8432, 8432, 8432, 8432, 8432, 8431, 8431, 8431, 
    8431, 8431, 8431, 8678, 8402, 8402, 8402, 8402, 8402, 8402,
  8669, 8779, 8427, 8427, 8426, 8426, 8427, 8427, 8427, 8426, 8426, 8426, 
    8426, 8426, 8426, 8677, 8424, 8424, 8424, 8424, 8424, 8424,
  8632, 8752, 8379, 8381, 8382, 8384, 8386, 8387, 8387, 8389, 8389, 8389, 
    8389, 8389, 8389, 8707, 8478, 8478, 8478, 8478, 8477, 8478,
  8858, 8970, 8381, 8382, 8383, 8384, 8385, 8386, 8386, 8387, 8387, 8387, 
    8387, 8387, 8387, 8778, 8436, 8436, 8436, 8436, 8435, 8436,
  8838, 8948, 8419, 8417, 8416, 8415, 8415, 8414, 8413, 8411, 8411, 8411, 
    8411, 8411, 8411, 8744, 8348, 8348, 8348, 8348, 8348, 8348,
  8839, 8949, 8596, 8593, 8591, 8589, 8588, 8587, 8586, 8582, 8582, 8582, 
    8582, 8582, 8582, 8820, 8474, 8474, 8474, 8474, 8474, 8474,
  8797, 8905, 8726, 8720, 8716, 8712, 8710, 8708, 8706, 8699, 8699, 8699, 
    8699, 8699, 8699, 8820, 8480, 8480, 8480, 8480, 8480, 8480,
  8872, 8974, 8794, 8788, 8783, 8780, 8778, 8776, 8774, 8767, 8767, 8767, 
    8767, 8767, 8767, 8868, 8556, 8556, 8556, 8556, 8556, 8556,
  8910, 9020, 8779, 8775, 8771, 8769, 8768, 8766, 8764, 8759, 8759, 8759, 
    8759, 8759, 8759, 8934, 8595, 8595, 8595, 8595, 8595, 8595,
  8887, 9000, 8741, 8740, 8739, 8738, 8738, 8738, 8737, 8736, 8736, 8736, 
    8736, 8736, 8736, 8950, 8694, 8694, 8694, 8694, 8694, 8694,
  8865, 8982, 8719, 8718, 8717, 8716, 8717, 8716, 8716, 8714, 8714, 8714, 
    8714, 8714, 8714, 8948, 8678, 8678, 8678, 8678, 8678, 8678,
  8832, 8945, 8700, 8696, 8694, 8692, 8691, 8690, 8689, 8685, 8685, 8685, 
    8685, 8685, 8685, 8879, 8565, 8565, 8565, 8565, 8565, 8565,
  8874, 8985, 8729, 8725, 8723, 8720, 8719, 8718, 8716, 8712, 8712, 8712, 
    8712, 8712, 8712, 8903, 8572, 8572, 8572, 8572, 8572, 8572,
  8870, 8978, 8771, 8772, 8773, 8774, 8775, 8776, 8776, 8778, 8778, 8778, 
    8778, 8778, 8778, 8957, 8836, 8836, 8836, 8836, 8836, 8836,
  8859, 8970, 8764, 8767, 8769, 8770, 8773, 8774, 8775, 8778, 8778, 8778, 
    8778, 8778, 8778, 8984, 8894, 8894, 8894, 8894, 8894, 8894,
  8757, 8877, 8674, 8680, 8684, 8686, 8690, 8692, 8694, 8700, 8700, 8700, 
    8700, 8700, 8700, 8950, 8913, 8913, 8913, 8913, 8913, 8913,
  8634, 8758, 8551, 8562, 8569, 8575, 8582, 8585, 8589, 8601, 8601, 8601, 
    8601, 8601, 8601, 8901, 9006, 9006, 9006, 9006, 9006, 9006,
  8327, 8472, 8189, 8204, 8215, 8223, 8232, 8237, 8242, 8259, 8259, 8259, 
    8259, 8259, 8259, 8707, 8828, 8828, 8828, 8828, 8828, 8828,
  8071, 8231, 7851, 7867, 7877, 7886, 7895, 7900, 7905, 7923, 7923, 7923, 
    7923, 7923, 7923, 8481, 8506, 8506, 8506, 8506, 8506, 8506,
  7730, 7907, 7570, 7586, 7598, 7607, 7616, 7622, 7628, 7646, 7646, 7646, 
    7646, 7646, 7646, 8256, 8274, 8274, 8274, 8274, 8274, 8274,
  7079, 7289, 6923, 6952, 6973, 6989, 7006, 7016, 7026, 7060, 7060, 7060, 
    7060, 7060, 7060, 7886, 8180, 8180, 8180, 8180, 8180, 8180,
  6820, 7046, 6524, 6554, 6574, 6590, 6606, 6617, 6627, 6660, 6660, 6660, 
    6660, 6660, 6660, 7625, 7766, 7766, 7766, 7766, 7766, 7766,
  6464, 6685, 6537, 6564, 6583, 6597, 6611, 6621, 6631, 6662, 6662, 6662, 
    6662, 6662, 6662, 7680, 7800, 7927, 7927, 7927, 7927, 7927,
  6562, 6823, 6206, 6245, 6273, 6294, 6315, 6329, 6343, 6386, 6386, 6386, 
    6386, 6386, 6386, 7602, 7857, 7857, 7857, 7857, 7857, 7857,
  6425, 6676, 6777, 6806, 6827, 6843, 6858, 6868, 6879, 6912, 6912, 6912, 
    6912, 6912, 6912, 7738, 8045, 8165, 8165, 8165, 8165, 8165,
  6765, 6997, 7126, 7152, 7170, 7184, 7198, 7206, 7216, 7245, 7245, 7245, 
    7245, 7245, 7245, 7936, 8233, 8342, 8342, 8342, 8342, 8342,
  6977, 7186, 7324, 7347, 7363, 7375, 7387, 7395, 7404, 7429, 7429, 7429, 
    7429, 7429, 7429, 8018, 8308, 8410, 8410, 8410, 8410, 8410,
  7176, 7370, 7410, 7430, 7445, 7456, 7466, 7473, 7482, 7505, 7505, 7505, 
    7505, 7505, 7505, 8133, 8327, 8426, 8426, 8426, 8426, 8426,
  7372, 7554, 7501, 7519, 7533, 7543, 7553, 7559, 7567, 7589, 7589, 7589, 
    7589, 7589, 7589, 8264, 8365, 8463, 8463, 8463, 8463, 8463,
  7430, 7589, 7389, 7406, 7418, 7427, 7436, 7441, 7449, 7468, 7468, 7468, 
    7468, 7468, 7468, 8236, 8228, 8329, 8329, 8329, 8329, 8329,
  7459, 7611, 7467, 7482, 7494, 7503, 7511, 7516, 7523, 7541, 7541, 7541, 
    7541, 7541, 7541, 8220, 8253, 8349, 8349, 8349, 8349, 8349,
  7471, 7649, 7636, 7654, 7667, 7677, 7686, 7692, 7700, 7720, 7720, 7720, 
    7720, 7720, 7720, 8321, 8444, 8537, 8537, 8537, 8537, 8537,
  7372, 7569, 7582, 7602, 7616, 7627, 7638, 7644, 7652, 7675, 7675, 7675, 
    7675, 7675, 7675, 8315, 8458, 8554, 8554, 8554, 8554, 8554,
  7273, 7475, 7463, 7484, 7499, 7511, 7522, 7529, 7537, 7561, 7561, 7561, 
    7561, 7561, 7561, 8260, 8396, 8496, 8496, 8496, 8496, 8496,
  7241, 7440, 7313, 7334, 7349, 7361, 7372, 7379, 7388, 7412, 7412, 7412, 
    7412, 7412, 7412, 8236, 8284, 8388, 8388, 8388, 8388, 8388,
  7133, 7342, 7282, 7304, 7321, 7333, 7344, 7352, 7361, 7387, 7387, 7387, 
    7387, 7387, 7387, 8177, 8286, 8391, 8391, 8391, 8391, 8391,
  7014, 7235, 7266, 7289, 7307, 7319, 7332, 7340, 7349, 7376, 7376, 7376, 
    7376, 7376, 7376, 8114, 8305, 8410, 8410, 8410, 8410, 8410,
  6767, 6997, 7077, 7103, 7121, 7135, 7148, 7157, 7167, 7196, 7196, 7196, 
    7196, 7196, 7196, 7937, 8193, 8303, 8303, 8303, 8303, 8303,
  6519, 6775, 6797, 6826, 6847, 6863, 6878, 6888, 6900, 6933, 6933, 6933, 
    6933, 6933, 6933, 7846, 8071, 8192, 8192, 8192, 8192, 8192,
  6281, 6528, 6297, 6328, 6349, 6366, 6382, 6392, 6404, 6439, 6439, 6439, 
    6439, 6439, 6439, 7650, 7707, 7842, 7842, 7842, 7842, 7842,
  6061, 6293, 6035, 6065, 6086, 6102, 6118, 6128, 6140, 6175, 6175, 6175, 
    6175, 6175, 6175, 7406, 7480, 7620, 7620, 7620, 7620, 7620,
  6008, 6237, 6013, 6042, 6063, 6080, 6095, 6105, 6117, 6151, 6151, 6151, 
    6151, 6151, 6151, 7341, 7452, 7593, 7593, 7593, 7593, 7593,
  6491, 6662, 6334, 6384, 6419, 6445, 6471, 6488, 6506, 6561, 6561, 6561, 
    6561, 6561, 6561, 7513, 8409, 8409, 8409, 8409, 8409, 8409,
  6825, 6991, 6693, 6731, 6758, 6778, 6797, 6810, 6824, 6866, 6866, 6866, 
    6866, 6866, 6866, 7641, 8274, 8274, 8274, 8274, 8274, 8274,
  7276, 7489, 7409, 7437, 7456, 7471, 7485, 7494, 7504, 7535, 7535, 7535, 
    7535, 7535, 7535, 8113, 8564, 8564, 8564, 8564, 8564, 8564,
  7417, 7569, 7582, 7597, 7609, 7617, 7625, 7630, 7637, 7654, 7654, 7654, 
    7654, 7654, 7654, 8161, 8329, 8421, 8421, 8421, 8421, 8421,
  7712, 7853, 7841, 7854, 7864, 7871, 7878, 7883, 7889, 7904, 7904, 7904, 
    7904, 7904, 7904, 8369, 8486, 8570, 8570, 8570, 8570, 8570,
  7925, 8065, 8084, 8096, 8105, 8112, 8118, 8122, 8128, 8141, 8141, 8141, 
    8141, 8141, 8141, 8539, 8655, 8733, 8733, 8733, 8733, 8733,
  7965, 8088, 8095, 8105, 8113, 8119, 8124, 8127, 8132, 8144, 8144, 8144, 
    8144, 8144, 8144, 8503, 8615, 8691, 8691, 8691, 8691, 8691,
  7995, 8101, 8100, 8109, 8115, 8120, 8125, 8127, 8132, 8141, 8141, 8141, 
    8141, 8141, 8141, 8455, 8569, 8644, 8644, 8644, 8644, 8644,
  8108, 8321, 8386, 8380, 8376, 8372, 8369, 8366, 8363, 8356, 8356, 8356, 
    8356, 8356, 8356, 8397, 8111, 8111, 8111, 8111, 8111, 8111,
  8115, 8312, 8359, 8351, 8346, 8341, 8337, 8333, 8330, 8321, 8321, 8321, 
    8321, 8321, 8321, 8309, 8006, 8006, 8006, 8006, 8006, 8006,
  8221, 8411, 8479, 8466, 8458, 8451, 8444, 8439, 8435, 8421, 8421, 8421, 
    8421, 8421, 8421, 8316, 7949, 7949, 7949, 7949, 7949, 7949,
  8183, 8409, 8599, 8583, 8571, 8562, 8554, 8547, 8541, 8523, 8523, 8523, 
    8523, 8523, 8523, 8358, 7901, 7901, 7901, 7901, 7901, 7901,
  8070, 8332, 8589, 8572, 8560, 8551, 8543, 8536, 8530, 8511, 8511, 8511, 
    8511, 8511, 8511, 8385, 7879, 7879, 7879, 7879, 7879, 7879,
  7778, 8090, 8464, 8448, 8437, 8428, 8419, 8413, 8407, 8389, 8389, 8389, 
    8389, 8389, 8389, 8295, 7776, 7776, 7776, 7776, 7776, 7776,
  7749, 8081, 8492, 8475, 8464, 8455, 8446, 8440, 8434, 8415, 8415, 8415, 
    8415, 8415, 8415, 8338, 7783, 7783, 7783, 7783, 7783, 7784,
  8782, 8899, 8984, 8983, 8983, 8983, 8984, 8983, 8983, 8983, 8983, 8983, 
    8983, 8983, 8983, 9041, 8979, 8979, 8979, 8979, 8979, 8979,
  8910, 9014, 9115, 9110, 9106, 9104, 9102, 9100, 9098, 9093, 9093, 9093, 
    9093, 9093, 9093, 9063, 8916, 8916, 8916, 8916, 8916, 8916,
  8811, 8918, 8951, 8949, 8949, 8948, 8948, 8948, 8947, 8946, 8946, 8946, 
    8946, 8946, 8946, 8981, 8913, 8913, 8913, 8913, 8913, 8913,
  8972, 9068, 9060, 9055, 9051, 9048, 9047, 9045, 9043, 9038, 9038, 9038, 
    9038, 9038, 9038, 9031, 8862, 8862, 8862, 8862, 8862, 8862,
  8873, 8969, 9009, 9004, 9001, 8998, 8997, 8995, 8993, 8988, 8988, 8988, 
    8988, 8988, 8988, 8956, 8818, 8818, 8818, 8818, 8818, 8818,
  9043, 9132, 9036, 9030, 9026, 9022, 9020, 9018, 9016, 9009, 9009, 9009, 
    9009, 9009, 9009, 9009, 8792, 8792, 8792, 8792, 8792, 8792,
  9260, 9324, 9187, 9173, 9163, 9156, 9150, 9145, 9140, 9125, 9125, 9125, 
    9125, 9125, 9125, 9000, 8622, 8622, 8622, 8622, 8622, 8622,
  9047, 9141, 8975, 8975, 8975, 8974, 8975, 8975, 8975, 8974, 8974, 8974, 
    8974, 8974, 8974, 9067, 8964, 8964, 8964, 8964, 8964, 8964,
  8957, 9057, 8929, 8930, 8931, 8931, 8933, 8933, 8934, 8935, 8935, 8935, 
    8935, 8935, 8935, 9047, 8991, 8991, 8991, 8991, 8991, 8991,
  8944, 9045, 8916, 8916, 8916, 8917, 8918, 8918, 8918, 8919, 8919, 8919, 
    8919, 8919, 8919, 9027, 8946, 8946, 8946, 8946, 8946, 8946,
  8819, 8920, 8736, 8733, 8732, 8730, 8730, 8729, 8728, 8725, 8725, 8725, 
    8725, 8725, 8725, 8837, 8640, 8640, 8640, 8640, 8640, 8640,
  8308, 8441, 8285, 8289, 8291, 8293, 8296, 8298, 8299, 8303, 8303, 8303, 
    8303, 8303, 8303, 8562, 8446, 8446, 8446, 8446, 8446, 8446,
  8643, 8756, 8514, 8514, 8515, 8515, 8517, 8517, 8517, 8518, 8518, 8518, 
    8518, 8518, 8518, 8730, 8560, 8560, 8560, 8560, 8560, 8560,
  8904, 8999, 8734, 8727, 8721, 8717, 8714, 8712, 8709, 8700, 8700, 8700, 
    8700, 8700, 8700, 8799, 8426, 8426, 8426, 8426, 8426, 8426,
  9031, 9124, 8912, 8907, 8903, 8900, 8898, 8897, 8895, 8889, 8889, 8889, 
    8889, 8889, 8889, 8975, 8708, 8708, 8708, 8708, 8708, 8708,
  8894, 9004, 8707, 8708, 8708, 8708, 8710, 8710, 8710, 8711, 8711, 8711, 
    8711, 8711, 8711, 8942, 8744, 8744, 8744, 8744, 8744, 8744,
  8838, 8948, 8639, 8640, 8641, 8642, 8643, 8643, 8644, 8645, 8645, 8645, 
    8645, 8645, 8645, 8886, 8693, 8693, 8693, 8693, 8693, 8693,
  9074, 9167, 8784, 8783, 8782, 8781, 8782, 8781, 8781, 8779, 8779, 8779, 
    8779, 8779, 8779, 8978, 8742, 8742, 8742, 8742, 8742, 8742,
  9107, 9197, 8840, 8838, 8836, 8835, 8835, 8834, 8833, 8831, 8831, 8831, 
    8831, 8831, 8831, 8998, 8757, 8757, 8757, 8757, 8757, 8757,
  9072, 9165, 8847, 8846, 8844, 8843, 8843, 8843, 8842, 8840, 8840, 8840, 
    8840, 8840, 8840, 9000, 8785, 8785, 8785, 8785, 8785, 8785,
  8988, 9085, 8811, 8809, 8808, 8808, 8808, 8807, 8807, 8805, 8805, 8805, 
    8805, 8805, 8805, 8962, 8759, 8759, 8759, 8759, 8759, 8759,
  8829, 8933, 8520, 8521, 8521, 8521, 8522, 8523, 8523, 8523, 8523, 8523, 
    8523, 8523, 8523, 8785, 8552, 8552, 8552, 8552, 8552, 8552,
  8349, 8476, 8139, 8143, 8146, 8148, 8152, 8153, 8155, 8159, 8159, 8159, 
    8159, 8159, 8159, 8494, 8324, 8324, 8324, 8324, 8324, 8324,
  8823, 8929, 8601, 8602, 8602, 8602, 8604, 8604, 8604, 8604, 8604, 8604, 
    8604, 8604, 8604, 8832, 8634, 8634, 8634, 8634, 8634, 8634,
  8773, 8896, 8645, 8651, 8655, 8658, 8662, 8664, 8666, 8672, 8672, 8672, 
    8672, 8672, 8672, 8969, 8896, 8896, 8896, 8896, 8896, 8896,
  8795, 8911, 8704, 8707, 8708, 8710, 8712, 8713, 8714, 8717, 8717, 8717, 
    8717, 8717, 8717, 8941, 8822, 8822, 8822, 8822, 8822, 8822,
  8887, 8987, 8642, 8642, 8642, 8642, 8643, 8643, 8643, 8643, 8643, 8643, 
    8643, 8643, 8643, 8852, 8647, 8647, 8647, 8647, 8647, 8647,
  8989, 9085, 8679, 8678, 8677, 8676, 8677, 8676, 8676, 8674, 8674, 8674, 
    8674, 8674, 8674, 8892, 8634, 8634, 8634, 8634, 8634, 8634,
  8930, 9043, 8681, 8687, 8691, 8694, 8698, 8700, 8702, 8708, 8708, 8708, 
    8708, 8708, 8708, 9025, 8936, 8936, 8936, 8936, 8936, 8936,
  8976, 9092, 8764, 8772, 8778, 8782, 8788, 8790, 8793, 8803, 8803, 8803, 
    8803, 8803, 8803, 9129, 9123, 9123, 9123, 9123, 9123, 9123,
  8935, 9052, 8702, 8709, 8714, 8718, 8723, 8725, 8727, 8735, 8735, 8735, 
    8735, 8735, 8735, 9065, 9004, 9004, 9004, 9004, 9004, 9004,
  8966, 9082, 8748, 8756, 8762, 8767, 8772, 8775, 8778, 8788, 8788, 8788, 
    8788, 8788, 8788, 9115, 9119, 9119, 9119, 9119, 9119, 9119,
  8954, 9065, 8675, 8680, 8684, 8687, 8691, 8692, 8694, 8700, 8700, 8700, 
    8700, 8700, 8700, 9013, 8905, 8905, 8905, 8905, 8905, 8905,
  8987, 9095, 8755, 8758, 8761, 8763, 8766, 8767, 8768, 8772, 8772, 8772, 
    8772, 8772, 8772, 9041, 8915, 8915, 8915, 8915, 8915, 8915,
  8985, 9092, 8726, 8729, 8731, 8732, 8735, 8736, 8737, 8740, 8740, 8740, 
    8740, 8740, 8740, 9011, 8852, 8852, 8852, 8852, 8852, 8852,
  8954, 9056, 8664, 8663, 8663, 8662, 8663, 8662, 8662, 8661, 8661, 8661, 
    8661, 8661, 8661, 8902, 8635, 8635, 8635, 8635, 8635, 8635,
  8920, 9023, 8669, 8666, 8663, 8662, 8661, 8660, 8659, 8656, 8656, 8656, 
    8656, 8656, 8656, 8866, 8555, 8555, 8555, 8555, 8555, 8555,
  8917, 9023, 8588, 8590, 8591, 8592, 8594, 8594, 8595, 8597, 8597, 8597, 
    8597, 8597, 8597, 8890, 8668, 8668, 8668, 8668, 8668, 8668,
  8915, 9017, 8660, 8656, 8654, 8652, 8651, 8650, 8648, 8644, 8644, 8644, 
    8644, 8644, 8644, 8849, 8517, 8517, 8517, 8517, 8517, 8517,
  8865, 8964, 8612, 8609, 8607, 8606, 8605, 8605, 8604, 8601, 8601, 8601, 
    8601, 8601, 8601, 8794, 8513, 8513, 8513, 8513, 8513, 8513,
  8950, 9047, 8654, 8652, 8650, 8649, 8649, 8648, 8648, 8645, 8645, 8645, 
    8645, 8645, 8645, 8855, 8578, 8578, 8578, 8578, 8578, 8578,
  8929, 9031, 8725, 8723, 8722, 8721, 8721, 8720, 8720, 8718, 8718, 8718, 
    8718, 8718, 8718, 8909, 8659, 8659, 8659, 8659, 8659, 8659,
  8920, 9021, 8647, 8645, 8643, 8642, 8641, 8641, 8640, 8637, 8637, 8637, 
    8637, 8637, 8637, 8851, 8554, 8554, 8554, 8554, 8554, 8554,
  9007, 9103, 8751, 8745, 8740, 8736, 8734, 8732, 8729, 8722, 8722, 8722, 
    8722, 8722, 8722, 8881, 8481, 8481, 8481, 8481, 8481, 8481,
  8975, 9073, 8880, 8871, 8866, 8861, 8858, 8855, 8852, 8843, 8843, 8843, 
    8843, 8843, 8843, 8921, 8547, 8547, 8547, 8547, 8547, 8547,
  8865, 8971, 8884, 8883, 8882, 8881, 8881, 8880, 8880, 8878, 8878, 8878, 
    8878, 8878, 8878, 8971, 8827, 8827, 8826, 8826, 8826, 8826,
  8839, 8947, 8791, 8790, 8790, 8789, 8790, 8790, 8789, 8788, 8788, 8788, 
    8788, 8788, 8788, 8927, 8766, 8766, 8766, 8766, 8766, 8766,
  8876, 8983, 8722, 8720, 8718, 8717, 8717, 8716, 8715, 8713, 8713, 8713, 
    8713, 8713, 8713, 8898, 8643, 8643, 8643, 8643, 8643, 8643,
  8928, 9032, 8639, 8631, 8626, 8622, 8619, 8616, 8614, 8605, 8605, 8605, 
    8605, 8605, 8605, 8812, 8332, 8332, 8332, 8332, 8332, 8332,
  8793, 8901, 8544, 8543, 8542, 8542, 8542, 8542, 8541, 8540, 8540, 8540, 
    8540, 8540, 8540, 8785, 8512, 8512, 8512, 8512, 8512, 8512,
  8895, 8998, 8799, 8792, 8787, 8784, 8782, 8779, 8777, 8770, 8770, 8770, 
    8770, 8770, 8770, 8879, 8537, 8537, 8537, 8537, 8537, 8537,
  8856, 8964, 8807, 8807, 8807, 8807, 8808, 8808, 8808, 8808, 8808, 8808, 
    8808, 8808, 8808, 8956, 8822, 8822, 8822, 8822, 8822, 8822,
  8996, 9102, 8853, 8855, 8856, 8858, 8860, 8860, 8861, 8864, 8864, 8864, 
    8864, 8864, 8864, 9070, 8955, 8955, 8955, 8955, 8955, 8955,
  9047, 9158, 8888, 8897, 8904, 8909, 8914, 8917, 8921, 8931, 8931, 8931, 
    8931, 8931, 8931, 9211, 9281, 9281, 9281, 9281, 9281, 9281,
  8900, 9018, 8721, 8734, 8742, 8749, 8757, 8761, 8766, 8780, 8780, 8780, 
    8780, 8780, 8780, 9125, 9263, 9263, 9263, 9263, 9263, 9263,
  8674, 8803, 8555, 8566, 8574, 8579, 8586, 8590, 8594, 8606, 8606, 8606, 
    8606, 8606, 8606, 8952, 9019, 9019, 9019, 9019, 9019, 9019,
  8376, 8519, 8255, 8270, 8281, 8288, 8297, 8302, 8307, 8324, 8324, 8324, 
    8324, 8324, 8324, 8753, 8884, 8884, 8884, 8884, 8884, 8884,
  8054, 8212, 7919, 7935, 7947, 7955, 7965, 7970, 7976, 7994, 7994, 7994, 
    7994, 7994, 7994, 8505, 8609, 8609, 8609, 8609, 8609, 8609,
  7635, 7817, 7510, 7533, 7549, 7562, 7575, 7583, 7591, 7617, 7617, 7617, 
    7617, 7617, 7617, 8269, 8496, 8496, 8496, 8496, 8496, 8496,
  7209, 7409, 6979, 7006, 7024, 7039, 7054, 7064, 7073, 7103, 7103, 7103, 
    7103, 7103, 7103, 7908, 8122, 8122, 8122, 8122, 8122, 8122,
  6750, 6975, 6909, 6934, 6953, 6967, 6980, 6989, 6999, 7029, 7029, 7029, 
    7029, 7029, 7029, 7928, 8077, 8194, 8194, 8194, 8194, 8194,
  6558, 6750, 6464, 6488, 6506, 6519, 6531, 6540, 6549, 6577, 6577, 6577, 
    6577, 6577, 6577, 7659, 7674, 7801, 7801, 7801, 7801, 7801,
  6509, 6733, 6684, 6711, 6730, 6744, 6758, 6767, 6778, 6808, 6808, 6808, 
    6808, 6808, 6808, 7716, 7912, 8034, 8034, 8034, 8034, 8034,
  6669, 6904, 7068, 7094, 7113, 7127, 7141, 7150, 7161, 7190, 7190, 7190, 
    7190, 7190, 7190, 7869, 8206, 8317, 8317, 8317, 8317, 8317,
  6950, 7175, 7317, 7341, 7358, 7371, 7384, 7392, 7402, 7429, 7429, 7429, 
    7429, 7429, 7429, 8061, 8348, 8451, 8451, 8451, 8451, 8451,
  7171, 7380, 7438, 7460, 7476, 7487, 7499, 7506, 7515, 7540, 7540, 7540, 
    7540, 7540, 7540, 8194, 8393, 8493, 8493, 8493, 8493, 8493,
  7333, 7512, 7427, 7446, 7460, 7470, 7480, 7486, 7494, 7515, 7515, 7515, 
    7515, 7515, 7515, 8222, 8310, 8410, 8410, 8410, 8410, 8410,
  7460, 7626, 7493, 7510, 7523, 7532, 7541, 7547, 7554, 7573, 7573, 7573, 
    7573, 7573, 7573, 8278, 8315, 8412, 8412, 8412, 8412, 8412,
  7526, 7671, 7453, 7468, 7479, 7488, 7496, 7501, 7507, 7525, 7525, 7525, 
    7525, 7525, 7525, 8261, 8236, 8334, 8334, 8334, 8334, 8334,
  7532, 7690, 7586, 7602, 7614, 7622, 7631, 7636, 7643, 7661, 7661, 7661, 
    7661, 7661, 7661, 8304, 8358, 8452, 8452, 8452, 8452, 8452,
  7416, 7608, 7590, 7610, 7624, 7634, 7645, 7651, 7659, 7681, 7681, 7681, 
    7681, 7681, 7681, 8338, 8457, 8553, 8553, 8553, 8553, 8553,
  7299, 7506, 7499, 7521, 7536, 7548, 7559, 7566, 7575, 7599, 7599, 7599, 
    7599, 7599, 7599, 8301, 8433, 8532, 8532, 8532, 8532, 8532,
  7233, 7443, 7310, 7332, 7348, 7360, 7372, 7380, 7389, 7414, 7414, 7414, 
    7414, 7414, 7414, 8279, 8316, 8421, 8421, 8421, 8421, 8421,
  7157, 7352, 7118, 7139, 7155, 7166, 7178, 7185, 7194, 7219, 7219, 7219, 
    7219, 7219, 7219, 8165, 8138, 8248, 8248, 8248, 8248, 8248,
  7116, 7310, 7150, 7172, 7187, 7199, 7210, 7217, 7226, 7251, 7251, 7251, 
    7251, 7251, 7251, 8118, 8157, 8265, 8265, 8265, 8265, 8265,
  7058, 7278, 7259, 7282, 7300, 7312, 7325, 7333, 7342, 7369, 7369, 7369, 
    7369, 7369, 7369, 8157, 8300, 8406, 8406, 8406, 8406, 8406,
  6957, 7187, 7267, 7291, 7309, 7322, 7335, 7344, 7354, 7381, 7381, 7381, 
    7381, 7381, 7381, 8095, 8326, 8431, 8431, 8431, 8431, 8431,
  6783, 7033, 7008, 7036, 7056, 7071, 7085, 7095, 7106, 7137, 7137, 7137, 
    7137, 7137, 7137, 8050, 8204, 8319, 8319, 8319, 8319, 8319,
  6584, 6835, 6773, 6802, 6823, 6838, 6853, 6863, 6874, 6907, 6907, 6907, 
    6907, 6907, 6907, 7897, 8047, 8168, 8168, 8168, 8168, 8168,
  6478, 6730, 6649, 6678, 6699, 6715, 6730, 6740, 6752, 6786, 6786, 6786, 
    6786, 6786, 6786, 7813, 7961, 8086, 8086, 8086, 8086, 8086,
  6457, 6693, 6718, 6746, 6765, 6780, 6795, 6804, 6815, 6847, 6847, 6847, 
    6847, 6847, 6847, 7715, 7962, 8083, 8083, 8083, 8083, 8083,
  6760, 6987, 6874, 6910, 6935, 6954, 6972, 6984, 6997, 7036, 7036, 7036, 
    7036, 7036, 7036, 7777, 8358, 8358, 8358, 8358, 8358, 8358,
  7112, 7300, 7185, 7220, 7245, 7263, 7281, 7293, 7306, 7345, 7345, 7345, 
    7345, 7345, 7345, 7959, 8648, 8648, 8648, 8648, 8648, 8648,
  7425, 7697, 7714, 7736, 7751, 7761, 7772, 7779, 7787, 7810, 7810, 7810, 
    7810, 7810, 7810, 8393, 8588, 8587, 8588, 8588, 8588, 8588,
  7480, 7637, 7665, 7680, 7692, 7700, 7709, 7714, 7721, 7738, 7738, 7738, 
    7738, 7738, 7738, 8234, 8405, 8495, 8495, 8495, 8495, 8495,
  7748, 7876, 7792, 7804, 7813, 7820, 7826, 7830, 7835, 7849, 7849, 7849, 
    7849, 7849, 7849, 8354, 8414, 8499, 8499, 8499, 8499, 8499,
  7887, 8009, 7952, 7963, 7971, 7977, 7983, 7986, 7991, 8003, 8003, 8003, 
    8003, 8003, 8003, 8438, 8510, 8591, 8591, 8591, 8591, 8591,
  7994, 8114, 8099, 8109, 8116, 8122, 8127, 8130, 8135, 8146, 8146, 8146, 
    8146, 8146, 8146, 8515, 8607, 8684, 8684, 8684, 8684, 8684,
  8099, 8224, 8247, 8257, 8264, 8270, 8275, 8278, 8283, 8294, 8294, 8294, 
    8294, 8294, 8294, 8619, 8726, 8799, 8799, 8799, 8799, 8799,
  8138, 8347, 8379, 8374, 8370, 8367, 8365, 8362, 8360, 8355, 8355, 8355, 
    8355, 8355, 8355, 8436, 8156, 8156, 8156, 8156, 8156, 8156,
  8227, 8432, 8531, 8521, 8514, 8509, 8504, 8500, 8496, 8485, 8485, 8485, 
    8485, 8485, 8485, 8426, 8109, 8109, 8109, 8109, 8109, 8109,
  8350, 8557, 8649, 8635, 8625, 8618, 8611, 8605, 8600, 8585, 8585, 8585, 
    8585, 8585, 8585, 8493, 8059, 8059, 8059, 8059, 8059, 8060,
  8360, 8576, 8694, 8677, 8665, 8656, 8647, 8641, 8635, 8616, 8616, 8616, 
    8616, 8616, 8616, 8494, 7976, 7976, 7976, 7976, 7976, 7976,
  8235, 8506, 8751, 8732, 8719, 8708, 8698, 8691, 8684, 8663, 8663, 8663, 
    8663, 8663, 8663, 8551, 7946, 7945, 7945, 7945, 7946, 7946,
  7969, 8301, 8708, 8687, 8673, 8662, 8651, 8644, 8636, 8613, 8613, 8613, 
    8613, 8613, 8613, 8502, 7840, 7839, 7839, 7839, 7840, 7840,
  7822, 8188, 8706, 8682, 8665, 8652, 8640, 8631, 8622, 8596, 8596, 8596, 
    8596, 8596, 8596, 8432, 7696, 7696, 7696, 7696, 7696, 7696,
  8759, 8871, 8999, 8997, 8996, 8995, 8995, 8995, 8994, 8992, 8992, 8992, 
    8992, 8992, 8992, 8999, 8938, 8938, 8938, 8938, 8938, 8938,
  8608, 8729, 8903, 8903, 8902, 8902, 8902, 8902, 8902, 8901, 8901, 8901, 
    8901, 8901, 8901, 8924, 8887, 8887, 8887, 8887, 8887, 8887,
  8793, 8898, 8986, 8983, 8981, 8980, 8980, 8979, 8978, 8975, 8975, 8975, 
    8975, 8975, 8975, 8968, 8894, 8894, 8894, 8894, 8894, 8894,
  9039, 9124, 9144, 9135, 9129, 9125, 9122, 9119, 9116, 9107, 9107, 9107, 
    9107, 9107, 9107, 9019, 8808, 8808, 8808, 8808, 8808, 8808,
  8877, 8975, 8975, 8970, 8968, 8965, 8964, 8963, 8961, 8956, 8956, 8956, 
    8956, 8956, 8956, 8954, 8810, 8810, 8810, 8810, 8810, 8810,
  9234, 9306, 9244, 9230, 9221, 9214, 9207, 9203, 9198, 9183, 9183, 9183, 
    9183, 9183, 9183, 9054, 8692, 8692, 8692, 8692, 8692, 8692,
  9084, 9163, 8891, 8885, 8881, 8877, 8875, 8873, 8870, 8863, 8863, 8863, 
    8863, 8863, 8863, 8913, 8638, 8638, 8638, 8638, 8638, 8638,
  9012, 9109, 8979, 8979, 8980, 8980, 8981, 8981, 8981, 8981, 8981, 8981, 
    8981, 8981, 8981, 9073, 9003, 9003, 9003, 9003, 9003, 9003,
  8945, 9047, 8918, 8920, 8920, 8921, 8922, 8923, 8923, 8925, 8925, 8925, 
    8925, 8925, 8925, 9037, 8977, 8977, 8977, 8977, 8977, 8977,
  8886, 8978, 8798, 8792, 8789, 8786, 8785, 8783, 8781, 8775, 8775, 8775, 
    8775, 8775, 8775, 8837, 8597, 8597, 8597, 8597, 8597, 8597,
  8909, 9001, 8841, 8837, 8834, 8832, 8831, 8829, 8828, 8823, 8823, 8823, 
    8823, 8823, 8823, 8881, 8675, 8676, 8676, 8676, 8676, 8676,
  8717, 8817, 8683, 8678, 8675, 8673, 8672, 8670, 8669, 8664, 8664, 8664, 
    8664, 8664, 8664, 8733, 8511, 8511, 8511, 8511, 8511, 8511,
  8760, 8864, 8659, 8658, 8657, 8657, 8657, 8657, 8656, 8655, 8655, 8655, 
    8655, 8655, 8655, 8801, 8633, 8633, 8633, 8633, 8633, 8633,
  9042, 9134, 8981, 8971, 8964, 8959, 8954, 8951, 8947, 8936, 8936, 8936, 
    8936, 8936, 8936, 8960, 8572, 8572, 8572, 8572, 8572, 8572,
  9037, 9130, 8903, 8898, 8894, 8891, 8889, 8887, 8885, 8878, 8878, 8878, 
    8878, 8878, 8878, 8969, 8679, 8679, 8679, 8679, 8679, 8679,
  8900, 9004, 8710, 8710, 8710, 8709, 8710, 8710, 8710, 8710, 8710, 8710, 
    8710, 8710, 8710, 8916, 8714, 8714, 8714, 8714, 8714, 8714,
  9023, 9117, 8728, 8728, 8727, 8727, 8728, 8728, 8727, 8727, 8727, 8727, 
    8727, 8727, 8727, 8935, 8715, 8715, 8715, 8715, 8715, 8715,
  9110, 9195, 8855, 8852, 8850, 8848, 8848, 8847, 8845, 8842, 8842, 8842, 
    8842, 8842, 8842, 8971, 8734, 8734, 8734, 8734, 8734, 8734,
  9141, 9227, 8863, 8860, 8857, 8856, 8855, 8854, 8853, 8849, 8849, 8849, 
    8849, 8849, 8849, 8999, 8745, 8745, 8745, 8745, 8745, 8745,
  9136, 9222, 8826, 8824, 8823, 8823, 8823, 8822, 8822, 8820, 8820, 8820, 
    8820, 8820, 8820, 8997, 8778, 8778, 8778, 8778, 8778, 8778,
  8796, 8899, 8491, 8492, 8493, 8493, 8495, 8495, 8495, 8496, 8496, 8496, 
    8496, 8496, 8496, 8757, 8539, 8539, 8539, 8539, 8539, 8539,
  8735, 8843, 8500, 8502, 8503, 8504, 8505, 8506, 8506, 8508, 8508, 8508, 
    8508, 8508, 8508, 8754, 8571, 8571, 8571, 8571, 8571, 8571,
  8842, 8948, 8587, 8588, 8589, 8589, 8591, 8591, 8591, 8592, 8592, 8592, 
    8592, 8592, 8592, 8840, 8634, 8634, 8634, 8634, 8634, 8634,
  8778, 8886, 8576, 8576, 8575, 8575, 8576, 8576, 8575, 8575, 8575, 8575, 
    8575, 8575, 8575, 8796, 8566, 8566, 8566, 8566, 8566, 8566,
  8756, 8868, 8528, 8528, 8529, 8529, 8531, 8531, 8531, 8531, 8531, 8531, 
    8531, 8531, 8531, 8791, 8563, 8563, 8563, 8563, 8563, 8563,
  8807, 8919, 8507, 8508, 8509, 8510, 8512, 8513, 8513, 8515, 8515, 8515, 
    8515, 8515, 8515, 8818, 8584, 8584, 8584, 8584, 8584, 8584,
  8822, 8937, 8597, 8601, 8604, 8606, 8610, 8611, 8613, 8618, 8618, 8618, 
    8618, 8618, 8618, 8920, 8790, 8790, 8790, 8790, 8790, 8790,
  8930, 9031, 8585, 8583, 8583, 8582, 8582, 8582, 8581, 8580, 8580, 8580, 
    8580, 8580, 8580, 8842, 8545, 8545, 8545, 8545, 8545, 8545,
  8891, 9007, 8565, 8573, 8578, 8582, 8587, 8589, 8592, 8600, 8600, 8600, 
    8600, 8600, 8600, 8977, 8885, 8885, 8885, 8885, 8885, 8885,
  8767, 8889, 8448, 8457, 8463, 8467, 8473, 8476, 8479, 8488, 8488, 8488, 
    8488, 8488, 8488, 8892, 8821, 8821, 8821, 8821, 8821, 8821,
  8890, 9006, 8603, 8609, 8614, 8617, 8621, 8624, 8626, 8633, 8633, 8633, 
    8633, 8633, 8633, 8983, 8882, 8882, 8882, 8882, 8882, 8882,
  8936, 9049, 8627, 8633, 8637, 8641, 8645, 8647, 8649, 8655, 8655, 8655, 
    8655, 8655, 8655, 8997, 8883, 8883, 8883, 8883, 8883, 8883,
  9077, 9169, 8769, 8766, 8764, 8762, 8761, 8760, 8759, 8756, 8756, 8756, 
    8756, 8756, 8756, 8949, 8653, 8653, 8653, 8653, 8652, 8653,
  9108, 9197, 8856, 8854, 8852, 8851, 8851, 8850, 8849, 8847, 8847, 8847, 
    8847, 8847, 8847, 9001, 8773, 8773, 8773, 8773, 8773, 8773,
  9184, 9271, 8912, 8906, 8903, 8900, 8898, 8896, 8894, 8888, 8888, 8888, 
    8888, 8888, 8888, 9029, 8701, 8701, 8701, 8701, 8701, 8701,
  9077, 9169, 8856, 8853, 8851, 8849, 8849, 8848, 8847, 8843, 8843, 8843, 
    8843, 8843, 8843, 8990, 8739, 8739, 8739, 8739, 8739, 8739,
  9110, 9204, 8882, 8879, 8877, 8875, 8875, 8874, 8873, 8869, 8869, 8869, 
    8869, 8869, 8869, 9031, 8764, 8764, 8764, 8764, 8764, 8764,
  9099, 9192, 8884, 8881, 8879, 8878, 8877, 8876, 8875, 8872, 8872, 8872, 
    8872, 8872, 8872, 9023, 8778, 8778, 8778, 8778, 8778, 8778,
  9040, 9134, 8825, 8822, 8820, 8818, 8818, 8816, 8815, 8812, 8812, 8812, 
    8812, 8812, 8812, 8965, 8711, 8711, 8711, 8711, 8711, 8711,
  9109, 9203, 9066, 9059, 9055, 9052, 9049, 9047, 9045, 9038, 9038, 9038, 
    9038, 9038, 9038, 9085, 8818, 8818, 8818, 8818, 8818, 8818,
  9042, 9138, 8785, 8783, 8781, 8780, 8780, 8779, 8778, 8776, 8776, 8776, 
    8776, 8776, 8776, 8965, 8702, 8702, 8702, 8702, 8702, 8702,
  9130, 9217, 8960, 8953, 8947, 8944, 8941, 8938, 8936, 8928, 8928, 8928, 
    8928, 8928, 8928, 9003, 8669, 8669, 8669, 8669, 8669, 8669,
  8883, 8987, 8632, 8631, 8631, 8631, 8632, 8631, 8631, 8631, 8631, 8631, 
    8631, 8631, 8631, 8864, 8626, 8626, 8626, 8626, 8626, 8626,
  8342, 8482, 8293, 8298, 8301, 8304, 8307, 8309, 8311, 8316, 8316, 8316, 
    8316, 8316, 8316, 8636, 8505, 8505, 8505, 8505, 8505, 8505,
  8565, 8691, 8406, 8409, 8411, 8413, 8415, 8417, 8418, 8421, 8421, 8421, 
    8421, 8421, 8421, 8720, 8543, 8543, 8543, 8543, 8543, 8543,
  8644, 8763, 8448, 8450, 8451, 8452, 8454, 8455, 8456, 8458, 8458, 8458, 
    8458, 8458, 8458, 8742, 8538, 8538, 8538, 8538, 8538, 8538,
  8931, 9033, 8601, 8597, 8595, 8593, 8592, 8590, 8589, 8584, 8584, 8584, 
    8584, 8584, 8584, 8825, 8447, 8447, 8447, 8447, 8447, 8447,
  8776, 8886, 8470, 8467, 8466, 8465, 8465, 8464, 8463, 8460, 8460, 8460, 
    8460, 8460, 8460, 8735, 8387, 8387, 8387, 8387, 8387, 8387,
  8908, 9017, 8649, 8641, 8635, 8631, 8627, 8625, 8621, 8612, 8612, 8612, 
    8612, 8612, 8612, 8827, 8310, 8310, 8310, 8310, 8310, 8310,
  8928, 9037, 8674, 8670, 8668, 8666, 8665, 8664, 8662, 8658, 8658, 8658, 
    8658, 8658, 8658, 8898, 8536, 8536, 8536, 8536, 8536, 8536,
  8867, 8979, 8697, 8696, 8695, 8694, 8694, 8694, 8693, 8692, 8692, 8692, 
    8692, 8692, 8692, 8916, 8651, 8651, 8651, 8651, 8651, 8651,
  8881, 8992, 8802, 8805, 8807, 8809, 8811, 8812, 8813, 8816, 8816, 8816, 
    8816, 8816, 8816, 9014, 8935, 8935, 8935, 8935, 8935, 8935,
  8983, 9093, 8891, 8897, 8901, 8904, 8908, 8910, 8912, 8919, 8919, 8919, 
    8919, 8919, 8919, 9139, 9145, 9145, 9145, 9145, 9145, 9145,
  8945, 9061, 8756, 8768, 8776, 8782, 8790, 8794, 8798, 8811, 8811, 8811, 
    8811, 8811, 8811, 9148, 9261, 9261, 9261, 9261, 9261, 9261,
  8936, 9044, 8756, 8759, 8760, 8761, 8763, 8764, 8765, 8767, 8767, 8767, 
    8767, 8767, 8767, 8998, 8858, 8858, 8858, 8858, 8858, 8858,
  8681, 8811, 8573, 8586, 8595, 8602, 8610, 8615, 8619, 8634, 8634, 8634, 
    8634, 8634, 8634, 8993, 9134, 9134, 9134, 9134, 9134, 9134,
  8308, 8454, 8343, 8358, 8370, 8378, 8387, 8393, 8399, 8416, 8416, 8416, 
    8416, 8416, 8416, 8789, 9020, 9020, 9020, 9020, 9020, 9020,
  7901, 8066, 7908, 7927, 7940, 7950, 7961, 7968, 7975, 7996, 7996, 7996, 
    7996, 7996, 7996, 8478, 8714, 8714, 8714, 8714, 8714, 8714,
  7662, 7840, 7461, 7479, 7492, 7502, 7513, 7519, 7526, 7546, 7546, 7546, 
    7546, 7546, 7546, 8186, 8247, 8247, 8247, 8247, 8247, 8247,
  7336, 7534, 6988, 7013, 7031, 7045, 7060, 7069, 7078, 7107, 7107, 7107, 
    7107, 7107, 7107, 7958, 8083, 8083, 8083, 8083, 8083, 8083,
  6837, 7022, 6788, 6810, 6826, 6838, 6849, 6857, 6866, 6891, 6891, 6891, 
    6891, 6891, 6891, 7855, 7881, 7999, 7999, 7999, 7999, 7999,
  6976, 7096, 6656, 6699, 6729, 6751, 6774, 6788, 6803, 6850, 6850, 6850, 
    6850, 6850, 6850, 7690, 8433, 8432, 8433, 8433, 8433, 8432,
  6738, 6953, 6863, 6888, 6906, 6919, 6932, 6941, 6951, 6979, 6979, 6979, 
    6979, 6979, 6979, 7880, 8018, 8135, 8135, 8135, 8135, 8135,
  6888, 7110, 7199, 7223, 7241, 7254, 7266, 7275, 7284, 7312, 7312, 7312, 
    7312, 7312, 7312, 8008, 8261, 8368, 8368, 8368, 8368, 8368,
  7156, 7365, 7449, 7471, 7487, 7499, 7510, 7518, 7527, 7551, 7551, 7551, 
    7551, 7551, 7551, 8177, 8401, 8501, 8501, 8501, 8501, 8501,
  7375, 7561, 7555, 7573, 7587, 7598, 7608, 7614, 7622, 7643, 7643, 7643, 
    7643, 7643, 7643, 8276, 8413, 8509, 8509, 8509, 8509, 8509,
  7523, 7668, 7482, 7497, 7508, 7517, 7525, 7529, 7536, 7553, 7553, 7553, 
    7553, 7553, 7553, 8255, 8256, 8353, 8353, 8353, 8353, 8353,
  7563, 7706, 7517, 7531, 7542, 7550, 7558, 7563, 7569, 7586, 7586, 7586, 
    7586, 7586, 7586, 8277, 8271, 8367, 8367, 8367, 8367, 8367,
  7541, 7678, 7469, 7483, 7494, 7502, 7509, 7514, 7520, 7537, 7537, 7537, 
    7537, 7537, 7537, 8242, 8226, 8323, 8323, 8323, 8323, 8323,
  7496, 7663, 7599, 7616, 7629, 7638, 7647, 7652, 7659, 7679, 7679, 7679, 
    7679, 7679, 7679, 8307, 8394, 8487, 8487, 8487, 8487, 8487,
  7350, 7547, 7529, 7549, 7564, 7575, 7585, 7592, 7600, 7623, 7623, 7623, 
    7623, 7623, 7623, 8302, 8426, 8524, 8524, 8524, 8524, 8524,
  7237, 7445, 7305, 7327, 7343, 7355, 7367, 7374, 7383, 7408, 7408, 7408, 
    7408, 7408, 7408, 8275, 8306, 8411, 8411, 8411, 8411, 8411,
  7147, 7340, 7031, 7052, 7068, 7080, 7091, 7098, 7107, 7132, 7132, 7132, 
    7132, 7132, 7132, 8157, 8075, 8189, 8189, 8189, 8189, 8189,
  7090, 7282, 6964, 6985, 7001, 7013, 7025, 7032, 7041, 7066, 7066, 7066, 
    7066, 7066, 7066, 8108, 8023, 8138, 8138, 8138, 8138, 8138,
  7094, 7299, 7084, 7107, 7123, 7135, 7147, 7155, 7164, 7190, 7190, 7190, 
    7190, 7190, 7190, 8151, 8141, 8252, 8252, 8252, 8252, 8252,
  7063, 7276, 7215, 7239, 7255, 7268, 7280, 7287, 7297, 7323, 7323, 7323, 
    7323, 7323, 7323, 8135, 8248, 8355, 8355, 8355, 8355, 8355,
  7030, 7249, 7244, 7267, 7285, 7297, 7310, 7318, 7327, 7354, 7354, 7354, 
    7354, 7354, 7354, 8129, 8289, 8395, 8395, 8395, 8395, 8395,
  7018, 7245, 7276, 7300, 7318, 7331, 7343, 7352, 7361, 7389, 7389, 7389, 
    7389, 7389, 7389, 8144, 8331, 8437, 8437, 8437, 8437, 8437,
  6925, 7155, 7102, 7127, 7146, 7159, 7172, 7181, 7191, 7220, 7220, 7220, 
    7220, 7220, 7220, 8088, 8216, 8327, 8327, 8327, 8327, 8327,
  6919, 7146, 7124, 7149, 7167, 7180, 7193, 7202, 7212, 7240, 7240, 7240, 
    7240, 7240, 7240, 8064, 8218, 8327, 8327, 8327, 8327, 8327,
  6823, 7046, 7108, 7133, 7151, 7164, 7177, 7185, 7195, 7223, 7223, 7223, 
    7223, 7223, 7223, 7959, 8197, 8306, 8306, 8306, 8306, 8306,
  7121, 7422, 7489, 7515, 7534, 7548, 7561, 7570, 7579, 7609, 7609, 7609, 
    7609, 7609, 7609, 8288, 8585, 8585, 8585, 8585, 8585, 8585,
  7242, 7471, 7426, 7452, 7470, 7484, 7497, 7505, 7514, 7543, 7543, 7543, 
    7543, 7543, 7543, 8105, 8493, 8492, 8492, 8492, 8493, 8492,
  7346, 7501, 7512, 7528, 7540, 7548, 7557, 7562, 7569, 7587, 7587, 7587, 
    7587, 7587, 7587, 8118, 8293, 8387, 8387, 8387, 8387, 8387,
  7583, 7735, 7750, 7764, 7775, 7783, 7791, 7796, 7802, 7819, 7819, 7819, 
    7819, 7819, 7819, 8302, 8451, 8538, 8538, 8538, 8538, 8538,
  7819, 7964, 7899, 7912, 7922, 7929, 7936, 7940, 7946, 7961, 7961, 7961, 
    7961, 7961, 7961, 8482, 8537, 8621, 8621, 8621, 8621, 8621,
  7931, 8053, 7996, 8006, 8014, 8020, 8026, 8029, 8034, 8046, 8046, 8046, 
    8046, 8046, 8046, 8477, 8541, 8621, 8621, 8621, 8621, 8621,
  8032, 8167, 8124, 8135, 8144, 8150, 8156, 8159, 8165, 8178, 8178, 8178, 
    8178, 8178, 8178, 8615, 8670, 8747, 8747, 8747, 8747, 8747,
  8104, 8227, 8187, 8197, 8204, 8210, 8215, 8218, 8223, 8234, 8234, 8234, 
    8234, 8234, 8234, 8625, 8682, 8757, 8757, 8757, 8757, 8757,
  8207, 8406, 8433, 8429, 8426, 8423, 8421, 8419, 8417, 8412, 8412, 8412, 
    8412, 8412, 8412, 8470, 8235, 8235, 8235, 8235, 8235, 8235,
  8223, 8405, 8432, 8425, 8420, 8416, 8412, 8409, 8407, 8399, 8399, 8399, 
    8399, 8399, 8399, 8372, 8124, 8124, 8124, 8124, 8124, 8124,
  8379, 8572, 8638, 8623, 8613, 8606, 8598, 8592, 8587, 8571, 8571, 8571, 
    8571, 8571, 8571, 8458, 8025, 8025, 8025, 8025, 8025, 8025,
  8436, 8632, 8684, 8669, 8659, 8652, 8644, 8638, 8633, 8617, 8617, 8617, 
    8617, 8617, 8617, 8530, 8066, 8066, 8066, 8066, 8066, 8066,
  8399, 8680, 8922, 8899, 8883, 8871, 8859, 8851, 8843, 8818, 8818, 8818, 
    8818, 8818, 8818, 8701, 7966, 7966, 7966, 7966, 7966, 7966,
  8080, 8390, 8707, 8689, 8677, 8667, 8658, 8652, 8645, 8625, 8625, 8625, 
    8625, 8625, 8625, 8576, 7961, 7961, 7961, 7961, 7961, 7961,
  7975, 8312, 8726, 8706, 8692, 8682, 8671, 8664, 8656, 8634, 8634, 8634, 
    8634, 8634, 8634, 8541, 7887, 7886, 7886, 7886, 7887, 7887,
  8778, 8891, 9027, 9025, 9024, 9023, 9023, 9023, 9022, 9021, 9021, 9021, 
    9021, 9021, 9021, 9033, 8975, 8974, 8974, 8974, 8974, 8974,
  8778, 8886, 8956, 8953, 8951, 8949, 8949, 8948, 8947, 8944, 8944, 8944, 
    8944, 8944, 8944, 8956, 8850, 8850, 8850, 8850, 8850, 8850,
  8880, 8980, 8908, 8906, 8905, 8904, 8904, 8903, 8903, 8901, 8901, 8901, 
    8901, 8901, 8901, 8960, 8847, 8847, 8847, 8847, 8847, 8847,
  8931, 9024, 8984, 8980, 8977, 8975, 8974, 8972, 8971, 8966, 8966, 8966, 
    8966, 8966, 8966, 8965, 8819, 8819, 8819, 8819, 8819, 8819,
  9278, 9343, 9301, 9285, 9273, 9265, 9257, 9251, 9245, 9227, 9227, 9227, 
    9227, 9227, 9227, 9042, 8627, 8627, 8627, 8627, 8627, 8627,
  8873, 8973, 8815, 8812, 8811, 8809, 8809, 8808, 8808, 8805, 8805, 8805, 
    8805, 8805, 8805, 8905, 8727, 8727, 8727, 8727, 8727, 8727,
  9020, 9117, 8946, 8946, 8946, 8946, 8947, 8947, 8947, 8947, 8947, 8947, 
    8947, 8947, 8947, 9059, 8956, 8956, 8956, 8956, 8956, 8956,
  8987, 9086, 8969, 8970, 8971, 8972, 8973, 8973, 8974, 8975, 8975, 8975, 
    8975, 8975, 8975, 9076, 9026, 9026, 9026, 9026, 9026, 9026,
  8975, 9074, 8960, 8960, 8960, 8960, 8961, 8961, 8961, 8961, 8961, 8961, 
    8961, 8961, 8961, 9051, 8975, 8975, 8975, 8975, 8975, 8975,
  9177, 9249, 9123, 9111, 9103, 9096, 9091, 9087, 9083, 9069, 9069, 9069, 
    9069, 9069, 9069, 8981, 8635, 8635, 8635, 8635, 8635, 8635,
  9007, 9096, 9015, 9005, 8997, 8991, 8987, 8983, 8979, 8967, 8967, 8967, 
    8967, 8967, 8967, 8933, 8581, 8581, 8581, 8581, 8581, 8581,
  8797, 8903, 8715, 8714, 8714, 8713, 8714, 8714, 8714, 8713, 8713, 8713, 
    8713, 8713, 8713, 8864, 8704, 8704, 8704, 8704, 8704, 8704,
  8861, 8963, 8750, 8748, 8747, 8746, 8746, 8746, 8745, 8743, 8743, 8743, 
    8743, 8743, 8743, 8882, 8685, 8685, 8685, 8685, 8685, 8685,
  8979, 9082, 8947, 8947, 8948, 8948, 8950, 8950, 8950, 8951, 8951, 8951, 
    8951, 8951, 8951, 9076, 8992, 8992, 8992, 8992, 8992, 8992,
  9100, 9195, 8953, 8946, 8942, 8938, 8936, 8934, 8932, 8924, 8924, 8924, 
    8924, 8924, 8924, 9028, 8698, 8698, 8698, 8698, 8698, 8698,
  9220, 9304, 9026, 9020, 9016, 9013, 9011, 9008, 9006, 9000, 9000, 9000, 
    9000, 9000, 9000, 9082, 8791, 8791, 8791, 8791, 8791, 8791,
  9135, 9222, 9014, 9009, 9005, 9002, 9000, 8998, 8997, 8991, 8991, 8991, 
    8991, 8991, 8991, 9051, 8805, 8805, 8805, 8805, 8805, 8805,
  9210, 9290, 8998, 8993, 8990, 8987, 8985, 8983, 8982, 8976, 8976, 8976, 
    8976, 8976, 8976, 9052, 8799, 8799, 8799, 8799, 8799, 8799,
  9232, 9313, 8876, 8873, 8870, 8868, 8867, 8866, 8865, 8861, 8861, 8861, 
    8861, 8861, 8861, 9027, 8742, 8742, 8742, 8742, 8742, 8742,
  8965, 9061, 8693, 8692, 8692, 8691, 8692, 8692, 8691, 8690, 8690, 8690, 
    8690, 8690, 8690, 8891, 8672, 8672, 8672, 8672, 8672, 8672,
  8928, 9028, 8704, 8704, 8704, 8704, 8705, 8705, 8705, 8705, 8705, 8705, 
    8705, 8705, 8705, 8904, 8709, 8709, 8709, 8709, 8709, 8709,
  9073, 9162, 8771, 8770, 8769, 8768, 8769, 8768, 8768, 8766, 8766, 8766, 
    8766, 8766, 8766, 8945, 8724, 8724, 8724, 8724, 8724, 8724,
  8808, 8913, 8604, 8605, 8605, 8605, 8606, 8606, 8606, 8607, 8607, 8607, 
    8607, 8607, 8607, 8822, 8627, 8627, 8627, 8627, 8627, 8627,
  8740, 8849, 8532, 8533, 8533, 8533, 8534, 8535, 8535, 8535, 8535, 8535, 
    8535, 8535, 8535, 8770, 8564, 8564, 8564, 8564, 8564, 8564,
  8764, 8877, 8469, 8470, 8471, 8472, 8473, 8474, 8474, 8476, 8476, 8476, 
    8476, 8476, 8476, 8778, 8534, 8534, 8534, 8534, 8534, 8534,
  8791, 8914, 8627, 8636, 8642, 8646, 8652, 8654, 8657, 8667, 8667, 8667, 
    8667, 8667, 8667, 8996, 8991, 8990, 8991, 8991, 8990, 8990,
  8879, 8980, 8601, 8600, 8600, 8600, 8601, 8600, 8600, 8600, 8600, 8600, 
    8600, 8600, 8600, 8826, 8594, 8594, 8594, 8594, 8594, 8594,
  8923, 9018, 8646, 8645, 8644, 8644, 8644, 8644, 8643, 8642, 8642, 8642, 
    8642, 8642, 8642, 8843, 8618, 8618, 8618, 8618, 8618, 8618,
  8783, 8903, 8463, 8470, 8476, 8479, 8484, 8487, 8489, 8497, 8497, 8497, 
    8497, 8497, 8497, 8887, 8780, 8780, 8780, 8780, 8780, 8780,
  8731, 8854, 8433, 8440, 8445, 8448, 8453, 8455, 8458, 8465, 8465, 8465, 
    8465, 8465, 8465, 8854, 8734, 8734, 8734, 8734, 8734, 8734,
  8819, 8937, 8549, 8554, 8557, 8560, 8563, 8565, 8567, 8572, 8572, 8572, 
    8572, 8572, 8572, 8912, 8765, 8765, 8765, 8765, 8765, 8765,
  8918, 9030, 8639, 8644, 8648, 8651, 8655, 8656, 8658, 8664, 8664, 8664, 
    8664, 8664, 8664, 8984, 8871, 8871, 8871, 8871, 8871, 8871,
  9036, 9138, 8823, 8825, 8826, 8826, 8828, 8829, 8829, 8831, 8831, 8831, 
    8831, 8831, 8831, 9046, 8891, 8891, 8891, 8891, 8891, 8891,
  9141, 9229, 8884, 8882, 8880, 8878, 8878, 8877, 8876, 8873, 8873, 8873, 
    8873, 8873, 8873, 9024, 8787, 8787, 8787, 8787, 8787, 8787,
  9208, 9294, 8897, 8894, 8892, 8890, 8889, 8888, 8887, 8884, 8884, 8884, 
    8884, 8884, 8884, 9048, 8780, 8780, 8781, 8781, 8780, 8780,
  9212, 9298, 8900, 8897, 8895, 8893, 8892, 8891, 8890, 8886, 8886, 8886, 
    8886, 8886, 8886, 9053, 8775, 8775, 8775, 8775, 8775, 8775,
  9272, 9359, 8991, 8987, 8985, 8983, 8983, 8981, 8980, 8977, 8977, 8977, 
    8977, 8977, 8977, 9131, 8862, 8862, 8862, 8862, 8862, 8862,
  9377, 9459, 9224, 9216, 9210, 9205, 9201, 9198, 9195, 9186, 9186, 9186, 
    9186, 9186, 9186, 9226, 8873, 8873, 8873, 8873, 8873, 8873,
  9362, 9442, 9223, 9214, 9209, 9204, 9201, 9198, 9195, 9186, 9186, 9186, 
    9186, 9186, 9186, 9212, 8887, 8887, 8887, 8887, 8887, 8887,
  9236, 9323, 9009, 9005, 9002, 9000, 8999, 8998, 8996, 8992, 8992, 8992, 
    8992, 8992, 8992, 9120, 8855, 8855, 8855, 8855, 8855, 8855,
  9145, 9236, 8813, 8809, 8807, 8805, 8805, 8803, 8802, 8798, 8798, 8798, 
    8798, 8798, 8798, 8994, 8684, 8684, 8684, 8684, 8684, 8684,
  8651, 8771, 8419, 8422, 8424, 8426, 8428, 8429, 8430, 8434, 8434, 8434, 
    8434, 8434, 8434, 8750, 8560, 8560, 8560, 8560, 8560, 8560,
  8302, 8448, 8179, 8185, 8190, 8193, 8198, 8200, 8202, 8210, 8210, 8210, 
    8210, 8210, 8210, 8600, 8462, 8462, 8462, 8462, 8462, 8462,
  8262, 8408, 8173, 8179, 8183, 8185, 8189, 8191, 8193, 8200, 8200, 8200, 
    8200, 8200, 8200, 8568, 8419, 8419, 8419, 8419, 8419, 8419,
  8797, 8903, 8622, 8623, 8623, 8624, 8625, 8625, 8625, 8626, 8626, 8626, 
    8626, 8626, 8626, 8832, 8661, 8661, 8661, 8661, 8661, 8661,
  8639, 8759, 8455, 8457, 8459, 8460, 8462, 8463, 8463, 8466, 8466, 8466, 
    8466, 8466, 8466, 8744, 8554, 8554, 8554, 8554, 8554, 8554,
  8509, 8634, 8247, 8248, 8249, 8250, 8252, 8252, 8253, 8254, 8254, 8254, 
    8254, 8254, 8254, 8591, 8320, 8320, 8320, 8320, 8320, 8320,
  8597, 8714, 8308, 8307, 8307, 8307, 8308, 8308, 8307, 8307, 8307, 8307, 
    8307, 8307, 8307, 8613, 8305, 8305, 8305, 8305, 8305, 8305,
  8643, 8758, 8527, 8528, 8529, 8529, 8531, 8531, 8531, 8532, 8532, 8532, 
    8532, 8532, 8532, 8751, 8578, 8578, 8578, 8578, 8578, 8578,
  8705, 8819, 8491, 8491, 8491, 8491, 8492, 8492, 8492, 8492, 8492, 8492, 
    8492, 8492, 8492, 8749, 8500, 8500, 8500, 8500, 8500, 8500,
  8756, 8870, 8597, 8598, 8599, 8600, 8602, 8602, 8603, 8605, 8605, 8605, 
    8605, 8605, 8605, 8847, 8669, 8669, 8669, 8669, 8669, 8669,
  8718, 8846, 8678, 8691, 8699, 8706, 8713, 8718, 8722, 8736, 8736, 8736, 
    8736, 8736, 8736, 9053, 9210, 9210, 9210, 9210, 9210, 9210,
  8785, 8908, 8820, 8828, 8834, 8838, 8843, 8846, 8849, 8858, 8858, 8858, 
    8858, 8858, 8858, 9084, 9169, 9169, 9169, 9169, 9169, 9169,
  8794, 8920, 8809, 8822, 8831, 8838, 8846, 8851, 8856, 8870, 8870, 8870, 
    8870, 8870, 8870, 9155, 9372, 9372, 9372, 9372, 9372, 9372,
  8728, 8856, 8688, 8700, 8709, 8715, 8722, 8726, 8731, 8744, 8744, 8744, 
    8744, 8744, 8744, 9052, 9203, 9203, 9203, 9203, 9203, 9203,
  8433, 8574, 8443, 8458, 8469, 8477, 8486, 8491, 8496, 8513, 8513, 8513, 
    8513, 8513, 8513, 8873, 9086, 9086, 9086, 9086, 9086, 9086,
  8103, 8262, 8149, 8169, 8184, 8195, 8207, 8214, 8221, 8244, 8244, 8244, 
    8244, 8244, 8244, 8698, 9025, 9025, 9025, 9025, 9025, 9025,
  7750, 7923, 7796, 7821, 7838, 7851, 7865, 7874, 7882, 7910, 7910, 7910, 
    7910, 7910, 7910, 8437, 8840, 8840, 8840, 8840, 8840, 8840,
  7504, 7690, 7209, 7238, 7258, 7273, 7289, 7300, 7310, 7342, 7342, 7342, 
    7342, 7342, 7342, 8132, 8428, 8428, 8428, 8428, 8428, 8428,
  7363, 7575, 6949, 6981, 7002, 7019, 7037, 7048, 7058, 7093, 7093, 7093, 
    7093, 7093, 7093, 8082, 8266, 8266, 8266, 8266, 8266, 8266,
  6869, 7063, 6971, 6993, 7009, 7021, 7033, 7041, 7050, 7075, 7075, 7075, 
    7075, 7075, 7075, 7898, 8030, 8143, 8143, 8143, 8143, 8143,
  6833, 7047, 7110, 7134, 7151, 7164, 7176, 7184, 7194, 7221, 7221, 7221, 
    7221, 7221, 7221, 7933, 8185, 8295, 8295, 8295, 8295, 8295,
  6862, 7078, 7141, 7165, 7183, 7195, 7208, 7216, 7226, 7253, 7253, 7253, 
    7253, 7253, 7253, 7962, 8204, 8312, 8312, 8312, 8312, 8312,
  7097, 7297, 7368, 7390, 7405, 7417, 7428, 7435, 7444, 7468, 7468, 7468, 
    7468, 7468, 7468, 8092, 8320, 8421, 8421, 8421, 8421, 8421,
  7312, 7500, 7551, 7570, 7584, 7594, 7605, 7611, 7619, 7641, 7641, 7641, 
    7641, 7641, 7641, 8219, 8411, 8506, 8506, 8506, 8506, 8506,
  7506, 7662, 7625, 7641, 7653, 7661, 7669, 7674, 7681, 7699, 7699, 7699, 
    7699, 7699, 7699, 8262, 8376, 8468, 8468, 8468, 8468, 8468,
  7618, 7759, 7644, 7658, 7668, 7676, 7683, 7688, 7694, 7710, 7710, 7710, 
    7710, 7710, 7710, 8305, 8351, 8442, 8442, 8442, 8442, 8442,
  7590, 7730, 7614, 7628, 7639, 7646, 7654, 7658, 7665, 7681, 7681, 7681, 
    7681, 7681, 7681, 8280, 8331, 8423, 8423, 8423, 8423, 8423,
  7592, 7729, 7528, 7542, 7553, 7560, 7568, 7572, 7579, 7595, 7595, 7595, 
    7595, 7595, 7595, 8281, 8267, 8362, 8362, 8362, 8362, 8362,
  7470, 7642, 7595, 7612, 7625, 7634, 7643, 7649, 7657, 7676, 7676, 7676, 
    7676, 7676, 7676, 8304, 8404, 8498, 8498, 8498, 8498, 8498,
  7289, 7490, 7406, 7427, 7442, 7454, 7465, 7472, 7480, 7504, 7504, 7504, 
    7504, 7504, 7504, 8279, 8356, 8458, 8458, 8458, 8458, 8458,
  7160, 7353, 7168, 7190, 7205, 7216, 7228, 7235, 7243, 7268, 7268, 7268, 
    7268, 7268, 7268, 8153, 8171, 8280, 8280, 8280, 8280, 8280,
  7062, 7239, 6829, 6850, 6865, 6876, 6887, 6894, 6903, 6927, 6927, 6927, 
    6927, 6927, 6927, 8032, 7890, 8008, 8008, 8008, 8008, 8008,
  6959, 7143, 6855, 6877, 6892, 6904, 6915, 6923, 6931, 6956, 6956, 6956, 
    6956, 6956, 6956, 7958, 7921, 8037, 8037, 8037, 8037, 8037,
  6979, 7173, 7031, 7052, 7068, 7080, 7092, 7099, 7108, 7133, 7133, 7133, 
    7133, 7133, 7133, 7995, 8068, 8179, 8179, 8179, 8179, 8179,
  7085, 7295, 7214, 7237, 7253, 7265, 7277, 7285, 7294, 7320, 7320, 7320, 
    7320, 7320, 7320, 8143, 8241, 8348, 8348, 8348, 8348, 8348,
  7125, 7332, 7355, 7377, 7393, 7405, 7416, 7424, 7433, 7458, 7458, 7458, 
    7458, 7458, 7458, 8150, 8331, 8433, 8433, 8433, 8433, 8433,
  7182, 7390, 7385, 7407, 7423, 7435, 7446, 7454, 7463, 7487, 7487, 7487, 
    7487, 7487, 7487, 8204, 8353, 8455, 8455, 8455, 8455, 8455,
  7185, 7394, 7388, 7410, 7426, 7438, 7449, 7457, 7466, 7491, 7491, 7491, 
    7491, 7491, 7491, 8213, 8357, 8459, 8459, 8459, 8459, 8459,
  7147, 7364, 7381, 7404, 7420, 7433, 7444, 7452, 7461, 7487, 7487, 7487, 
    7487, 7487, 7487, 8212, 8375, 8477, 8477, 8477, 8477, 8477,
  7157, 7364, 7409, 7430, 7446, 7458, 7469, 7476, 7485, 7509, 7509, 7509, 
    7509, 7509, 7509, 8169, 8361, 8461, 8461, 8461, 8461, 8461,
  7221, 7415, 7426, 7446, 7461, 7472, 7482, 7489, 7497, 7520, 7520, 7520, 
    7520, 7520, 7520, 8176, 8338, 8437, 8437, 8437, 8437, 8437,
  7359, 7537, 7535, 7554, 7567, 7577, 7587, 7592, 7600, 7621, 7621, 7621, 
    7621, 7621, 7621, 8227, 8374, 8470, 8470, 8470, 8470, 8470,
  7504, 7655, 7596, 7611, 7623, 7631, 7639, 7644, 7650, 7668, 7668, 7668, 
    7668, 7668, 7668, 8241, 8340, 8432, 8432, 8432, 8432, 8432,
  7682, 7840, 7794, 7809, 7820, 7828, 7836, 7841, 7848, 7865, 7865, 7865, 
    7865, 7865, 7865, 8422, 8503, 8591, 8591, 8591, 8591, 8591,
  7802, 7942, 7846, 7859, 7869, 7876, 7883, 7887, 7893, 7908, 7908, 7908, 
    7908, 7908, 7908, 8452, 8490, 8575, 8575, 8575, 8575, 8575,
  7890, 8017, 7942, 7953, 7962, 7968, 7974, 7977, 7983, 7996, 7996, 7996, 
    7996, 7996, 7996, 8465, 8517, 8598, 8598, 8598, 8598, 8598,
  7993, 8115, 8108, 8118, 8126, 8131, 8137, 8140, 8145, 8156, 8156, 8156, 
    8156, 8156, 8156, 8523, 8620, 8697, 8697, 8697, 8697, 8697,
  8123, 8254, 8310, 8320, 8328, 8333, 8339, 8342, 8347, 8358, 8358, 8358, 
    8358, 8358, 8358, 8658, 8784, 8856, 8856, 8856, 8856, 8856,
  8171, 8373, 8427, 8420, 8414, 8410, 8406, 8402, 8399, 8391, 8391, 8391, 
    8391, 8391, 8391, 8395, 8089, 8089, 8089, 8089, 8089, 8089,
  8341, 8534, 8596, 8582, 8573, 8565, 8558, 8553, 8548, 8533, 8533, 8533, 
    8533, 8533, 8533, 8434, 8021, 8021, 8021, 8021, 8021, 8021,
  8448, 8620, 8621, 8607, 8596, 8588, 8581, 8575, 8569, 8553, 8553, 8553, 
    8553, 8553, 8553, 8443, 7992, 7992, 7992, 7992, 7992, 7992,
  8579, 8781, 8864, 8845, 8831, 8821, 8811, 8804, 8796, 8775, 8775, 8775, 
    8775, 8775, 8775, 8620, 8049, 8049, 8049, 8049, 8049, 8049,
  8440, 8700, 8932, 8908, 8892, 8880, 8867, 8859, 8850, 8824, 8824, 8824, 
    8824, 8824, 8824, 8648, 7943, 7943, 7943, 7943, 7943, 7943,
  8177, 8492, 8840, 8819, 8805, 8794, 8783, 8775, 8768, 8745, 8745, 8745, 
    8745, 8745, 8745, 8643, 7969, 7969, 7969, 7969, 7969, 7969,
  8022, 8353, 8752, 8731, 8717, 8706, 8695, 8687, 8680, 8656, 8656, 8656, 
    8656, 8656, 8656, 8548, 7874, 7874, 7874, 7874, 7874, 7874,
  8737, 8851, 8943, 8942, 8941, 8940, 8940, 8940, 8939, 8938, 8938, 8938, 
    8938, 8938, 8938, 8972, 8893, 8893, 8893, 8893, 8893, 8893,
  8893, 8988, 8976, 8969, 8964, 8961, 8958, 8955, 8953, 8945, 8945, 8945, 
    8945, 8945, 8945, 8918, 8694, 8694, 8694, 8694, 8694, 8694,
  8957, 9045, 9087, 9081, 9077, 9074, 9072, 9070, 9068, 9061, 9061, 9061, 
    9061, 9061, 9061, 8988, 8856, 8856, 8856, 8856, 8856, 8856,
  9030, 9110, 9055, 9047, 9042, 9038, 9034, 9032, 9029, 9021, 9021, 9021, 
    9021, 9021, 9021, 8950, 8746, 8746, 8746, 8746, 8746, 8746,
  9041, 9127, 8959, 8953, 8949, 8946, 8945, 8943, 8941, 8935, 8935, 8935, 
    8935, 8935, 8935, 8963, 8744, 8744, 8744, 8744, 8744, 8744,
  9077, 9172, 9020, 9020, 9020, 9020, 9021, 9021, 9021, 9021, 9021, 9021, 
    9021, 9021, 9021, 9119, 9031, 9031, 9031, 9031, 9031, 9031,
  9023, 9120, 8971, 8971, 8971, 8971, 8972, 8972, 8972, 8972, 8972, 8972, 
    8972, 8972, 8972, 9077, 8987, 8987, 8987, 8987, 8987, 8987,
  8598, 8715, 8685, 8685, 8684, 8684, 8684, 8684, 8684, 8683, 8683, 8683, 
    8683, 8683, 8683, 8791, 8671, 8671, 8671, 8671, 8671, 8671,
  8921, 9013, 8891, 8886, 8883, 8881, 8879, 8878, 8876, 8871, 8871, 8871, 
    8871, 8871, 8871, 8907, 8711, 8711, 8711, 8711, 8712, 8711,
  9114, 9205, 9149, 9139, 9132, 9126, 9122, 9118, 9115, 9103, 9103, 9103, 
    9103, 9103, 9103, 9071, 8730, 8730, 8730, 8730, 8730, 8730,
  8884, 8986, 8833, 8831, 8829, 8827, 8827, 8826, 8825, 8822, 8822, 8822, 
    8822, 8822, 8822, 8924, 8731, 8731, 8731, 8731, 8731, 8731,
  8879, 8984, 8823, 8821, 8820, 8820, 8820, 8819, 8819, 8817, 8817, 8817, 
    8817, 8817, 8817, 8943, 8771, 8771, 8771, 8771, 8771, 8771,
  8847, 8950, 8797, 8794, 8792, 8790, 8790, 8788, 8787, 8784, 8784, 8784, 
    8784, 8784, 8784, 8887, 8676, 8676, 8676, 8676, 8676, 8676,
  9002, 9105, 8963, 8963, 8964, 8964, 8965, 8965, 8965, 8966, 8966, 8966, 
    8966, 8966, 8966, 9089, 8993, 8993, 8993, 8993, 8993, 8993,
  9018, 9122, 8976, 8977, 8977, 8978, 8979, 8980, 8980, 8981, 8981, 8981, 
    8981, 8981, 8981, 9120, 9032, 9032, 9032, 9032, 9032, 9032,
  9083, 9176, 8951, 8947, 8945, 8942, 8941, 8940, 8939, 8934, 8934, 8934, 
    8934, 8934, 8934, 9035, 8801, 8801, 8801, 8801, 8801, 8801,
  9097, 9184, 8855, 8852, 8850, 8848, 8848, 8847, 8845, 8842, 8842, 8842, 
    8842, 8842, 8842, 8978, 8740, 8740, 8740, 8740, 8740, 8740,
  9292, 9371, 9089, 9078, 9071, 9066, 9061, 9058, 9054, 9042, 9042, 9042, 
    9042, 9042, 9042, 9078, 8665, 8665, 8665, 8665, 8665, 8665,
  9165, 9249, 8857, 8854, 8852, 8851, 8850, 8849, 8848, 8844, 8844, 8844, 
    8844, 8844, 8844, 9000, 8741, 8741, 8741, 8741, 8741, 8741,
  8915, 9014, 8580, 8581, 8581, 8582, 8583, 8583, 8584, 8584, 8584, 8584, 
    8584, 8584, 8584, 8841, 8622, 8622, 8622, 8622, 8622, 8622,
  9112, 9198, 8793, 8792, 8790, 8789, 8790, 8789, 8788, 8786, 8786, 8786, 
    8786, 8786, 8786, 8965, 8733, 8733, 8733, 8733, 8733, 8733,
  9034, 9126, 8748, 8747, 8746, 8746, 8746, 8746, 8745, 8744, 8744, 8744, 
    8744, 8744, 8744, 8932, 8714, 8714, 8714, 8714, 8714, 8714,
  8846, 8950, 8584, 8585, 8585, 8585, 8586, 8586, 8587, 8587, 8587, 8587, 
    8587, 8587, 8587, 8825, 8612, 8612, 8612, 8612, 8612, 8612,
  8827, 8933, 8534, 8535, 8536, 8537, 8538, 8539, 8539, 8540, 8540, 8540, 
    8540, 8540, 8540, 8812, 8590, 8590, 8590, 8590, 8590, 8590,
  8826, 8933, 8513, 8513, 8513, 8513, 8513, 8514, 8513, 8513, 8513, 8513, 
    8513, 8513, 8513, 8790, 8521, 8521, 8521, 8521, 8521, 8521,
  8862, 8975, 8676, 8679, 8682, 8683, 8686, 8687, 8689, 8692, 8692, 8692, 
    8692, 8692, 8692, 8953, 8829, 8829, 8829, 8829, 8829, 8829,
  8724, 8828, 8434, 8434, 8434, 8434, 8435, 8435, 8435, 8435, 8435, 8435, 
    8435, 8435, 8435, 8683, 8449, 8449, 8449, 8449, 8449, 8449,
  8965, 9059, 8742, 8740, 8739, 8739, 8739, 8738, 8738, 8736, 8736, 8736, 
    8736, 8736, 8736, 8896, 8688, 8688, 8688, 8688, 8688, 8688,
  8862, 8981, 8655, 8662, 8668, 8671, 8676, 8679, 8681, 8689, 8689, 8689, 
    8689, 8689, 8689, 9015, 8971, 8971, 8971, 8971, 8971, 8971,
  8776, 8901, 8553, 8563, 8569, 8575, 8581, 8584, 8588, 8599, 8599, 8599, 
    8599, 8599, 8599, 8976, 8973, 8973, 8973, 8973, 8973, 8973,
  8762, 8883, 8456, 8463, 8467, 8471, 8475, 8477, 8480, 8487, 8487, 8487, 
    8487, 8487, 8487, 8864, 8739, 8739, 8739, 8739, 8739, 8739,
  8887, 8999, 8605, 8610, 8613, 8615, 8619, 8620, 8622, 8627, 8627, 8627, 
    8627, 8627, 8627, 8941, 8803, 8803, 8803, 8803, 8803, 8803,
  9022, 9123, 8742, 8743, 8743, 8744, 8745, 8745, 8746, 8746, 8746, 8746, 
    8746, 8746, 8746, 8991, 8783, 8783, 8783, 8783, 8783, 8783,
  9103, 9192, 8798, 8796, 8795, 8794, 8794, 8793, 8792, 8790, 8790, 8790, 
    8790, 8790, 8790, 8972, 8722, 8722, 8722, 8722, 8722, 8722,
  9209, 9292, 8939, 8936, 8934, 8932, 8931, 8930, 8929, 8925, 8925, 8925, 
    8925, 8925, 8925, 9060, 8818, 8818, 8818, 8818, 8818, 8818,
  9315, 9395, 8950, 8947, 8944, 8943, 8942, 8941, 8940, 8936, 8936, 8936, 
    8936, 8936, 8936, 9108, 8826, 8826, 8826, 8826, 8826, 8826,
  8799, 8911, 8520, 8522, 8523, 8524, 8526, 8527, 8528, 8529, 8529, 8529, 
    8529, 8529, 8529, 8827, 8606, 8606, 8606, 8606, 8606, 8606,
  8961, 9066, 8638, 8639, 8639, 8640, 8641, 8641, 8642, 8643, 8643, 8643, 
    8643, 8643, 8643, 8926, 8686, 8686, 8686, 8686, 8686, 8686,
  9336, 9419, 8944, 8941, 8939, 8937, 8936, 8935, 8933, 8929, 8929, 8929, 
    8929, 8929, 8929, 9127, 8808, 8808, 8808, 8808, 8808, 8808,
  9276, 9360, 8918, 8916, 8914, 8913, 8913, 8912, 8912, 8909, 8909, 8909, 
    8909, 8909, 8909, 9102, 8840, 8840, 8840, 8840, 8840, 8840,
  8912, 9019, 8518, 8519, 8521, 8521, 8523, 8524, 8524, 8526, 8526, 8526, 
    8526, 8526, 8526, 8855, 8596, 8596, 8596, 8596, 8596, 8596,
  8857, 8966, 8571, 8573, 8573, 8574, 8576, 8576, 8577, 8578, 8578, 8578, 
    8578, 8578, 8578, 8861, 8640, 8640, 8640, 8640, 8640, 8640,
  9136, 9225, 8868, 8865, 8863, 8861, 8861, 8860, 8859, 8855, 8855, 8855, 
    8855, 8855, 8855, 9014, 8753, 8753, 8753, 8753, 8753, 8753,
  8941, 9042, 8658, 8657, 8656, 8655, 8655, 8655, 8654, 8653, 8653, 8653, 
    8653, 8653, 8653, 8880, 8611, 8611, 8611, 8611, 8611, 8611,
  8848, 8955, 8712, 8707, 8704, 8702, 8700, 8699, 8697, 8692, 8692, 8692, 
    8692, 8692, 8692, 8849, 8529, 8529, 8529, 8529, 8529, 8529,
  8638, 8755, 8476, 8472, 8469, 8467, 8466, 8465, 8464, 8459, 8459, 8459, 
    8459, 8459, 8459, 8683, 8327, 8327, 8327, 8327, 8327, 8327,
  8696, 8820, 8554, 8551, 8550, 8549, 8549, 8548, 8547, 8545, 8545, 8545, 
    8545, 8545, 8545, 8804, 8480, 8480, 8480, 8480, 8480, 8480,
  8390, 8525, 8250, 8253, 8256, 8258, 8261, 8262, 8264, 8268, 8268, 8268, 
    8268, 8268, 8268, 8606, 8420, 8420, 8420, 8420, 8420, 8420,
  8389, 8529, 8221, 8235, 8244, 8251, 8259, 8264, 8268, 8283, 8283, 8283, 
    8283, 8283, 8283, 8715, 8792, 8792, 8792, 8792, 8792, 8792,
  8380, 8521, 8330, 8346, 8358, 8366, 8376, 8381, 8387, 8405, 8405, 8405, 
    8405, 8405, 8405, 8794, 9019, 9019, 9019, 9019, 9019, 9019,
  8371, 8513, 8363, 8378, 8388, 8395, 8404, 8409, 8414, 8430, 8430, 8430, 
    8430, 8430, 8430, 8796, 8973, 8973, 8973, 8973, 8973, 8973,
  8539, 8670, 8561, 8574, 8583, 8590, 8597, 8601, 8606, 8620, 8620, 8620, 
    8620, 8620, 8620, 8912, 9100, 9100, 9100, 9100, 9100, 9100,
  8476, 8613, 8533, 8541, 8546, 8550, 8555, 8558, 8561, 8569, 8569, 8569, 
    8569, 8569, 8569, 8837, 8863, 8863, 8863, 8863, 8863, 8863,
  8382, 8531, 8539, 8557, 8570, 8579, 8589, 8595, 8602, 8622, 8622, 8622, 
    8622, 8622, 8622, 8958, 9297, 9296, 9296, 9296, 9296, 9296,
  8206, 8363, 8381, 8402, 8416, 8427, 8438, 8445, 8453, 8476, 8476, 8476, 
    8476, 8476, 8476, 8851, 9247, 9247, 9247, 9247, 9247, 9247,
  8115, 8275, 8197, 8222, 8239, 8252, 8266, 8274, 8283, 8310, 8310, 8310, 
    8310, 8310, 8310, 8771, 9234, 9234, 9234, 9234, 9234, 9234,
  7826, 8000, 7741, 7768, 7786, 7800, 7815, 7824, 7834, 7863, 7863, 7863, 
    7863, 7863, 7863, 8478, 8856, 8856, 8856, 8856, 8856, 8856,
  7442, 7638, 7708, 7728, 7742, 7753, 7763, 7769, 7777, 7799, 7799, 7799, 
    7799, 7799, 7799, 8364, 8549, 8642, 8642, 8642, 8642, 8642,
  7310, 7511, 7378, 7399, 7415, 7426, 7437, 7444, 7453, 7477, 7477, 7477, 
    7477, 7477, 7477, 8304, 8340, 8444, 8444, 8444, 8444, 8444,
  7108, 7296, 7170, 7191, 7206, 7218, 7228, 7235, 7244, 7268, 7268, 7268, 
    7268, 7268, 7268, 8081, 8158, 8265, 8265, 8265, 8265, 8265,
  6917, 7116, 7190, 7212, 7228, 7240, 7251, 7259, 7268, 7293, 7293, 7293, 
    7293, 7293, 7293, 7936, 8189, 8295, 8295, 8295, 8295, 8295,
  6918, 7135, 7296, 7319, 7336, 7349, 7361, 7369, 7378, 7405, 7405, 7405, 
    7405, 7405, 7405, 7996, 8311, 8415, 8415, 8415, 8415, 8415,
  7045, 7251, 7374, 7396, 7412, 7424, 7436, 7443, 7452, 7477, 7477, 7477, 
    7477, 7477, 7477, 8064, 8339, 8440, 8440, 8440, 8440, 8440,
  7299, 7482, 7480, 7499, 7513, 7523, 7533, 7539, 7547, 7569, 7569, 7569, 
    7569, 7569, 7569, 8198, 8348, 8445, 8445, 8445, 8445, 8445,
  7490, 7662, 7634, 7652, 7664, 7673, 7683, 7688, 7696, 7715, 7715, 7715, 
    7715, 7715, 7715, 8316, 8434, 8528, 8528, 8528, 8528, 8528,
  7607, 7759, 7691, 7706, 7717, 7725, 7733, 7738, 7744, 7762, 7762, 7762, 
    7762, 7762, 7762, 8337, 8418, 8509, 8509, 8509, 8509, 8509,
  7699, 7843, 7795, 7808, 7818, 7826, 7833, 7837, 7843, 7859, 7859, 7859, 
    7859, 7859, 7859, 8371, 8459, 8546, 8546, 8546, 8546, 8546,
  7707, 7837, 7674, 7687, 7697, 7704, 7710, 7714, 7720, 7735, 7735, 7735, 
    7735, 7735, 7735, 8342, 8348, 8438, 8438, 8438, 8438, 8438,
  7604, 7734, 7596, 7609, 7619, 7626, 7633, 7637, 7643, 7658, 7658, 7658, 
    7658, 7658, 7658, 8249, 8286, 8377, 8377, 8377, 8377, 8377,
  7468, 7641, 7542, 7560, 7572, 7582, 7591, 7597, 7604, 7624, 7624, 7624, 
    7624, 7624, 7624, 8310, 8367, 8463, 8463, 8463, 8463, 8463,
  7324, 7508, 7405, 7425, 7439, 7449, 7459, 7465, 7474, 7496, 7496, 7496, 
    7496, 7496, 7496, 8236, 8302, 8402, 8402, 8402, 8402, 8402,
  7163, 7350, 7131, 7152, 7167, 7178, 7189, 7195, 7204, 7228, 7228, 7228, 
    7228, 7228, 7228, 8130, 8123, 8231, 8231, 8231, 8231, 8231,
  7026, 7204, 6985, 7005, 7020, 7031, 7042, 7048, 7057, 7081, 7081, 7081, 
    7081, 7081, 7081, 7979, 7994, 8105, 8105, 8105, 8105, 8105,
  6918, 7123, 6957, 6980, 6997, 7010, 7022, 7030, 7039, 7066, 7066, 7066, 
    7066, 7066, 7066, 7993, 8048, 8162, 8162, 8162, 8162, 8162,
  6972, 7179, 7068, 7091, 7108, 7120, 7132, 7140, 7149, 7176, 7176, 7176, 
    7176, 7176, 7176, 8043, 8133, 8244, 8244, 8244, 8244, 8244,
  7096, 7305, 7169, 7191, 7208, 7220, 7232, 7240, 7249, 7275, 7275, 7275, 
    7275, 7275, 7275, 8157, 8207, 8316, 8316, 8316, 8316, 8316,
  7237, 7444, 7364, 7386, 7401, 7413, 7425, 7432, 7441, 7465, 7465, 7465, 
    7465, 7465, 7465, 8257, 8337, 8440, 8440, 8440, 8440, 8440,
  7353, 7558, 7501, 7522, 7537, 7548, 7559, 7566, 7575, 7599, 7599, 7599, 
    7599, 7599, 7599, 8344, 8430, 8530, 8530, 8530, 8530, 8530,
  7370, 7566, 7554, 7574, 7588, 7599, 7609, 7616, 7624, 7647, 7647, 7647, 
    7647, 7647, 7647, 8314, 8441, 8538, 8538, 8538, 8538, 8538,
  7398, 7596, 7597, 7617, 7632, 7643, 7653, 7660, 7668, 7690, 7690, 7690, 
    7690, 7690, 7690, 8342, 8473, 8569, 8569, 8569, 8569, 8569,
  7421, 7613, 7618, 7638, 7652, 7662, 7673, 7679, 7687, 7709, 7709, 7709, 
    7709, 7709, 7709, 8340, 8473, 8568, 8568, 8568, 8568, 8568,
  7450, 7618, 7593, 7610, 7622, 7631, 7640, 7646, 7653, 7672, 7672, 7672, 
    7672, 7672, 7672, 8263, 8386, 8479, 8479, 8479, 8479, 8479,
  7528, 7686, 7597, 7613, 7625, 7633, 7642, 7647, 7654, 7672, 7672, 7672, 
    7672, 7672, 7672, 8295, 8361, 8454, 8454, 8454, 8454, 8454,
  7627, 7779, 7692, 7707, 7718, 7726, 7734, 7739, 7745, 7762, 7762, 7762, 
    7762, 7762, 7762, 8354, 8413, 8503, 8503, 8503, 8503, 8503,
  7693, 7832, 7734, 7747, 7757, 7765, 7772, 7776, 7782, 7797, 7797, 7797, 
    7797, 7797, 7797, 8352, 8403, 8490, 8490, 8490, 8490, 8490,
  7727, 7863, 7726, 7739, 7749, 7756, 7763, 7767, 7773, 7788, 7788, 7788, 
    7788, 7788, 7788, 8377, 8393, 8482, 8482, 8482, 8482, 8482,
  7857, 7994, 7969, 7981, 7991, 7997, 8004, 8007, 8013, 8027, 8027, 8027, 
    8027, 8027, 8027, 8473, 8564, 8645, 8645, 8645, 8645, 8645,
  7915, 8034, 8035, 8045, 8053, 8058, 8064, 8067, 8072, 8083, 8083, 8083, 
    8083, 8083, 8083, 8442, 8559, 8637, 8637, 8637, 8637, 8637,
  8051, 8164, 8241, 8249, 8256, 8261, 8266, 8268, 8273, 8283, 8283, 8283, 
    8283, 8283, 8283, 8521, 8687, 8759, 8759, 8759, 8759, 8759,
  8236, 8451, 8525, 8516, 8510, 8505, 8500, 8497, 8494, 8484, 8484, 8484, 
    8484, 8484, 8484, 8495, 8151, 8151, 8151, 8151, 8151, 8151,
  8359, 8553, 8639, 8623, 8612, 8603, 8595, 8588, 8582, 8564, 8564, 8564, 
    8564, 8564, 8564, 8415, 7951, 7951, 7951, 7951, 7951, 7951,
  8490, 8652, 8683, 8665, 8653, 8644, 8634, 8627, 8621, 8601, 8601, 8601, 
    8601, 8601, 8601, 8390, 7928, 7928, 7928, 7928, 7928, 7928,
  8620, 8820, 8939, 8913, 8896, 8883, 8869, 8860, 8851, 8823, 8823, 8823, 
    8823, 8823, 8823, 8559, 7877, 7877, 7877, 7877, 7877, 7877,
  8431, 8654, 8816, 8793, 8777, 8765, 8753, 8745, 8736, 8711, 8711, 8711, 
    8711, 8711, 8711, 8493, 7847, 7846, 7846, 7846, 7847, 7847,
  8176, 8472, 8827, 8803, 8786, 8773, 8761, 8752, 8743, 8716, 8716, 8716, 
    8716, 8716, 8716, 8506, 7809, 7809, 7809, 7809, 7809, 7809,
  8021, 8323, 8678, 8658, 8645, 8635, 8625, 8618, 8610, 8589, 8589, 8589, 
    8589, 8589, 8589, 8453, 7863, 7863, 7863, 7863, 7863, 7863,
  8789, 8892, 8948, 8942, 8937, 8934, 8932, 8930, 8928, 8921, 8921, 8921, 
    8921, 8921, 8921, 8900, 8708, 8708, 8708, 8708, 8708, 8708,
  8864, 8961, 9018, 9010, 9005, 9001, 8998, 8995, 8993, 8984, 8984, 8984, 
    8984, 8984, 8984, 8929, 8714, 8714, 8714, 8714, 8714, 8714,
  8971, 9063, 9005, 9001, 8998, 8996, 8995, 8994, 8992, 8988, 8988, 8988, 
    8988, 8988, 8988, 8994, 8854, 8854, 8854, 8854, 8854, 8854,
  9064, 9147, 8979, 8974, 8971, 8969, 8967, 8966, 8964, 8959, 8959, 8959, 
    8959, 8959, 8959, 8978, 8794, 8794, 8794, 8794, 8794, 8794,
  8577, 8698, 8665, 8666, 8667, 8667, 8669, 8669, 8669, 8670, 8670, 8670, 
    8670, 8670, 8670, 8807, 8717, 8717, 8717, 8717, 8717, 8717,
  9073, 9168, 9009, 9010, 9010, 9010, 9011, 9011, 9011, 9012, 9012, 9012, 
    9012, 9012, 9012, 9117, 9033, 9033, 9033, 9033, 9033, 9033,
  8945, 9039, 8907, 8903, 8901, 8899, 8897, 8896, 8895, 8890, 8890, 8890, 
    8890, 8890, 8890, 8943, 8753, 8753, 8753, 8753, 8753, 8753,
  9188, 9266, 9200, 9188, 9180, 9173, 9168, 9164, 9159, 9146, 9146, 9146, 
    9146, 9146, 9146, 9052, 8706, 8706, 8706, 8706, 8706, 8706,
  8983, 9077, 8944, 8939, 8936, 8933, 8931, 8929, 8927, 8922, 8922, 8922, 
    8922, 8922, 8922, 8968, 8741, 8741, 8741, 8741, 8741, 8741,
  8944, 9042, 8944, 8941, 8938, 8936, 8935, 8934, 8933, 8929, 8929, 8929, 
    8929, 8929, 8929, 8984, 8804, 8804, 8804, 8804, 8804, 8804,
  8966, 9070, 8986, 8981, 8978, 8975, 8974, 8972, 8970, 8965, 8965, 8965, 
    8965, 8965, 8965, 9035, 8798, 8798, 8798, 8798, 8798, 8798,
  8943, 9043, 8836, 8835, 8834, 8833, 8833, 8832, 8832, 8830, 8830, 8830, 
    8830, 8830, 8830, 8964, 8785, 8785, 8785, 8785, 8785, 8785,
  9061, 9162, 9037, 9028, 9021, 9017, 9013, 9010, 9006, 8996, 8996, 8996, 
    8996, 8996, 8996, 9050, 8670, 8670, 8670, 8670, 8670, 8670,
  8931, 9039, 8869, 8869, 8870, 8870, 8871, 8872, 8872, 8872, 8872, 8872, 
    8872, 8872, 8872, 9032, 8903, 8903, 8903, 8903, 8903, 8903,
  8958, 9064, 8867, 8865, 8864, 8863, 8863, 8863, 8862, 8860, 8860, 8860, 
    8860, 8860, 8860, 9016, 8809, 8809, 8809, 8809, 8809, 8809,
  9101, 9194, 9004, 9002, 8999, 8998, 8997, 8996, 8995, 8992, 8992, 8992, 
    8992, 8992, 8992, 9082, 8893, 8893, 8893, 8893, 8893, 8893,
  9188, 9272, 8979, 8973, 8968, 8965, 8962, 8960, 8958, 8950, 8950, 8950, 
    8950, 8950, 8950, 9032, 8717, 8717, 8717, 8717, 8717, 8717,
  9189, 9276, 9083, 9078, 9074, 9071, 9069, 9067, 9065, 9058, 9058, 9058, 
    9058, 9058, 9058, 9108, 8860, 8860, 8860, 8860, 8860, 8860,
  9123, 9210, 8815, 8811, 8809, 8807, 8806, 8805, 8804, 8800, 8800, 8800, 
    8800, 8800, 8800, 8967, 8685, 8685, 8685, 8685, 8685, 8685,
  9090, 9178, 8741, 8739, 8737, 8735, 8735, 8734, 8733, 8730, 8730, 8730, 
    8730, 8730, 8730, 8925, 8639, 8639, 8639, 8639, 8639, 8639,
  9071, 9162, 8741, 8737, 8735, 8733, 8731, 8730, 8729, 8724, 8724, 8724, 
    8724, 8724, 8724, 8918, 8586, 8586, 8586, 8586, 8586, 8586,
  8916, 9026, 8700, 8702, 8704, 8705, 8708, 8709, 8710, 8712, 8712, 8712, 
    8712, 8712, 8712, 8974, 8819, 8819, 8819, 8819, 8819, 8819,
  8902, 9005, 8579, 8577, 8576, 8575, 8575, 8575, 8574, 8572, 8572, 8572, 
    8572, 8572, 8572, 8824, 8520, 8520, 8520, 8520, 8520, 8520,
  8855, 8963, 8500, 8501, 8501, 8502, 8503, 8504, 8504, 8505, 8505, 8505, 
    8505, 8505, 8505, 8812, 8544, 8544, 8544, 8544, 8544, 8544,
  8914, 9024, 8721, 8724, 8726, 8728, 8730, 8731, 8732, 8736, 8736, 8736, 
    8736, 8736, 8736, 8988, 8857, 8857, 8857, 8857, 8857, 8857,
  8940, 9040, 8630, 8630, 8629, 8629, 8630, 8630, 8630, 8629, 8629, 8629, 
    8629, 8629, 8629, 8874, 8626, 8626, 8626, 8626, 8626, 8626,
  8900, 8999, 8564, 8563, 8562, 8561, 8562, 8562, 8561, 8560, 8560, 8560, 
    8560, 8560, 8560, 8804, 8534, 8534, 8534, 8534, 8534, 8534,
  8970, 9083, 8715, 8721, 8726, 8729, 8733, 8735, 8737, 8744, 8744, 8744, 
    8744, 8744, 8744, 9063, 8984, 8984, 8984, 8984, 8984, 8984,
  8858, 8976, 8590, 8599, 8605, 8609, 8615, 8618, 8621, 8631, 8631, 8631, 
    8631, 8631, 8631, 8996, 8969, 8969, 8969, 8969, 8969, 8969,
  8830, 8949, 8475, 8483, 8488, 8492, 8497, 8500, 8502, 8511, 8511, 8511, 
    8511, 8511, 8511, 8914, 8802, 8802, 8802, 8802, 8802, 8802,
  8845, 8961, 8443, 8450, 8454, 8458, 8462, 8465, 8467, 8474, 8474, 8474, 
    8474, 8474, 8474, 8882, 8726, 8726, 8726, 8726, 8726, 8726,
  8905, 9016, 8571, 8576, 8579, 8581, 8584, 8586, 8587, 8592, 8592, 8592, 
    8592, 8592, 8592, 8930, 8764, 8764, 8764, 8764, 8764, 8764,
  8985, 9089, 8718, 8719, 8719, 8720, 8721, 8721, 8721, 8722, 8722, 8722, 
    8722, 8722, 8722, 8968, 8755, 8755, 8755, 8755, 8755, 8755,
  9065, 9162, 8871, 8871, 8870, 8870, 8871, 8871, 8871, 8870, 8870, 8870, 
    8870, 8870, 8870, 9047, 8866, 8866, 8866, 8866, 8866, 8866,
  9240, 9326, 9020, 9017, 9015, 9013, 9013, 9012, 9011, 9007, 9007, 9007, 
    9007, 9007, 9007, 9133, 8906, 8906, 8906, 8906, 8906, 8906,
  9420, 9494, 9147, 9140, 9135, 9131, 9128, 9125, 9122, 9114, 9114, 9114, 
    9114, 9114, 9114, 9185, 8848, 8848, 8848, 8848, 8848, 8848,
  9349, 9430, 8980, 8977, 8975, 8974, 8973, 8972, 8971, 8968, 8968, 8968, 
    8968, 8968, 8968, 9146, 8874, 8874, 8874, 8874, 8874, 8874,
  9637, 9699, 9332, 9320, 9312, 9305, 9300, 9296, 9291, 9278, 9278, 9278, 
    9278, 9278, 9278, 9286, 8842, 8842, 8842, 8842, 8842, 8842,
  9599, 9666, 9300, 9289, 9281, 9275, 9270, 9266, 9262, 9250, 9250, 9250, 
    9250, 9250, 9250, 9282, 8844, 8844, 8844, 8844, 8844, 8844,
  9557, 9622, 9250, 9237, 9229, 9222, 9216, 9212, 9207, 9193, 9193, 9193, 
    9193, 9193, 9193, 9212, 8736, 8736, 8736, 8736, 8736, 8736,
  9261, 9344, 8969, 8966, 8964, 8962, 8961, 8960, 8959, 8955, 8955, 8955, 
    8955, 8955, 8955, 9101, 8845, 8845, 8845, 8845, 8845, 8845,
  9168, 9255, 9038, 9034, 9032, 9029, 9028, 9027, 9025, 9021, 9021, 9021, 
    9021, 9021, 9021, 9092, 8881, 8881, 8881, 8881, 8881, 8881,
  8970, 9068, 8748, 8745, 8743, 8741, 8741, 8740, 8738, 8735, 8735, 8735, 
    8735, 8735, 8735, 8911, 8637, 8637, 8637, 8637, 8637, 8637,
  8597, 8711, 8311, 8311, 8311, 8311, 8312, 8312, 8312, 8312, 8312, 8312, 
    8312, 8312, 8312, 8601, 8322, 8322, 8322, 8322, 8322, 8322,
  8653, 8775, 8428, 8428, 8427, 8427, 8428, 8428, 8427, 8427, 8427, 8427, 
    8427, 8427, 8427, 8725, 8417, 8417, 8417, 8417, 8417, 8417,
  8409, 8544, 8226, 8230, 8233, 8235, 8238, 8240, 8241, 8246, 8246, 8246, 
    8246, 8246, 8246, 8605, 8410, 8410, 8410, 8410, 8410, 8410,
  8281, 8424, 8061, 8071, 8078, 8084, 8090, 8094, 8097, 8108, 8108, 8108, 
    8108, 8108, 8108, 8561, 8498, 8498, 8498, 8498, 8498, 8498,
  8138, 8294, 7893, 7907, 7917, 7924, 7932, 7937, 7942, 7957, 7957, 7957, 
    7957, 7957, 7957, 8503, 8479, 8479, 8479, 8479, 8479, 8479,
  8097, 8251, 7965, 7980, 7991, 7999, 8009, 8014, 8020, 8037, 8037, 8037, 
    8037, 8037, 8037, 8523, 8627, 8627, 8627, 8627, 8627, 8627,
  8038, 8199, 8064, 8086, 8102, 8114, 8126, 8134, 8142, 8166, 8166, 8166, 
    8166, 8166, 8166, 8642, 9000, 9000, 9000, 9000, 9000, 9000,
  8095, 8257, 8228, 8253, 8271, 8284, 8298, 8307, 8316, 8345, 8345, 8345, 
    8345, 8345, 8345, 8794, 9302, 9302, 9302, 9302, 9302, 9302,
  8075, 8239, 8111, 8135, 8151, 8163, 8176, 8184, 8192, 8218, 8218, 8218, 
    8218, 8218, 8218, 8711, 9090, 9090, 9090, 9090, 9090, 9090,
  8026, 8189, 8028, 8050, 8065, 8076, 8088, 8096, 8103, 8127, 8127, 8127, 
    8127, 8127, 8127, 8624, 8933, 8933, 8933, 8933, 8933, 8933,
  7914, 8087, 7982, 8010, 8030, 8044, 8060, 8070, 8080, 8111, 8111, 8111, 
    8111, 8111, 8111, 8660, 9171, 9171, 9171, 9171, 9171, 9171,
  7876, 8071, 7961, 8000, 8028, 8049, 8071, 8085, 8099, 8143, 8143, 8143, 
    8143, 8143, 8143, 8857, 9630, 9630, 9630, 9630, 9630, 9630,
  7737, 7916, 7417, 7441, 7458, 7471, 7485, 7493, 7502, 7529, 7529, 7529, 
    7529, 7529, 7529, 8279, 8444, 8444, 8444, 8444, 8444, 8444,
  7670, 7852, 7317, 7339, 7354, 7366, 7378, 7386, 7393, 7418, 7418, 7418, 
    7418, 7418, 7418, 8182, 8244, 8244, 8244, 8244, 8244, 8244,
  7282, 7476, 7419, 7439, 7454, 7465, 7476, 7482, 7491, 7514, 7514, 7514, 
    7514, 7514, 7514, 8236, 8340, 8440, 8440, 8440, 8440, 8440,
  7119, 7313, 7208, 7229, 7244, 7256, 7267, 7274, 7283, 7307, 7307, 7307, 
    7307, 7307, 7307, 8113, 8203, 8310, 8310, 8310, 8310, 8310,
  7069, 7262, 7160, 7181, 7196, 7208, 7219, 7226, 7235, 7260, 7260, 7260, 
    7260, 7260, 7260, 8064, 8164, 8273, 8273, 8273, 8273, 8273,
  7065, 7270, 7322, 7344, 7360, 7372, 7383, 7391, 7400, 7425, 7425, 7425, 
    7425, 7425, 7425, 8087, 8303, 8406, 8406, 8406, 8406, 8406,
  7090, 7286, 7329, 7350, 7365, 7376, 7387, 7394, 7403, 7427, 7427, 7427, 
    7427, 7427, 7427, 8073, 8281, 8384, 8384, 8384, 8384, 8384,
  7240, 7413, 7367, 7385, 7399, 7409, 7419, 7425, 7433, 7454, 7454, 7454, 
    7454, 7454, 7454, 8115, 8245, 8344, 8344, 8344, 8344, 8344,
  7463, 7623, 7447, 7464, 7476, 7485, 7494, 7499, 7506, 7526, 7526, 7526, 
    7526, 7526, 7526, 8266, 8274, 8373, 8373, 8373, 8373, 8373,
  7600, 7757, 7718, 7734, 7745, 7753, 7761, 7766, 7773, 7791, 7791, 7791, 
    7791, 7791, 7791, 8347, 8448, 8538, 8538, 8538, 8538, 8538,
  7688, 7837, 7823, 7837, 7847, 7855, 7862, 7867, 7873, 7889, 7889, 7889, 
    7889, 7889, 7889, 8381, 8495, 8581, 8581, 8581, 8581, 8581,
  7751, 7891, 7824, 7837, 7847, 7854, 7861, 7865, 7871, 7887, 7887, 7887, 
    7887, 7887, 7887, 8409, 8484, 8571, 8571, 8571, 8571, 8571,
  7718, 7857, 7679, 7693, 7703, 7710, 7718, 7722, 7728, 7744, 7744, 7744, 
    7744, 7744, 7744, 8393, 8381, 8472, 8472, 8472, 8472, 8472,
  7649, 7804, 7700, 7715, 7727, 7735, 7743, 7748, 7754, 7772, 7772, 7772, 
    7772, 7772, 7772, 8390, 8432, 8523, 8523, 8523, 8523, 8523,
  7547, 7723, 7693, 7710, 7723, 7732, 7741, 7747, 7754, 7774, 7774, 7774, 
    7774, 7774, 7774, 8380, 8483, 8575, 8575, 8575, 8575, 8575,
  7342, 7534, 7441, 7461, 7475, 7486, 7497, 7503, 7512, 7534, 7534, 7534, 
    7534, 7534, 7534, 8287, 8354, 8455, 8455, 8455, 8455, 8455,
  7174, 7371, 7265, 7287, 7302, 7314, 7325, 7332, 7341, 7365, 7365, 7365, 
    7365, 7365, 7365, 8172, 8248, 8354, 8354, 8354, 8354, 8354,
  6992, 7203, 7056, 7080, 7097, 7109, 7122, 7130, 7139, 7166, 7166, 7166, 
    7166, 7166, 7166, 8081, 8137, 8249, 8249, 8249, 8249, 8249,
  6928, 7140, 7011, 7034, 7052, 7064, 7077, 7085, 7095, 7122, 7122, 7122, 
    7122, 7122, 7122, 8028, 8106, 8219, 8219, 8219, 8219, 8219,
  6966, 7175, 7028, 7052, 7069, 7081, 7094, 7102, 7111, 7138, 7138, 7138, 
    7138, 7138, 7138, 8052, 8113, 8225, 8225, 8225, 8225, 8225,
  7145, 7356, 7210, 7232, 7249, 7261, 7273, 7281, 7290, 7316, 7316, 7316, 
    7316, 7316, 7316, 8209, 8246, 8354, 8354, 8354, 8354, 8354,
  7359, 7546, 7384, 7404, 7418, 7429, 7439, 7446, 7454, 7476, 7476, 7476, 
    7476, 7476, 7476, 8288, 8299, 8401, 8401, 8401, 8401, 8401,
  7493, 7681, 7549, 7568, 7582, 7592, 7603, 7609, 7617, 7639, 7639, 7639, 
    7639, 7639, 7639, 8403, 8419, 8517, 8517, 8517, 8517, 8517,
  7514, 7708, 7600, 7620, 7634, 7644, 7655, 7661, 7669, 7691, 7691, 7691, 
    7691, 7691, 7691, 8439, 8470, 8566, 8566, 8566, 8566, 8566,
  7556, 7741, 7634, 7652, 7666, 7675, 7685, 7691, 7699, 7720, 7720, 7720, 
    7720, 7720, 7720, 8438, 8470, 8565, 8565, 8565, 8565, 8565,
  7594, 7777, 7658, 7676, 7690, 7699, 7709, 7715, 7722, 7743, 7743, 7743, 
    7743, 7743, 7743, 8464, 8481, 8575, 8575, 8575, 8575, 8575,
  7612, 7778, 7644, 7660, 7672, 7681, 7689, 7695, 7702, 7720, 7720, 7720, 
    7720, 7720, 7720, 8405, 8419, 8511, 8511, 8511, 8511, 8511,
  7624, 7780, 7648, 7663, 7675, 7683, 7691, 7696, 7703, 7721, 7721, 7721, 
    7721, 7721, 7721, 8378, 8397, 8489, 8489, 8489, 8489, 8489,
  7671, 7829, 7727, 7742, 7753, 7762, 7770, 7775, 7781, 7799, 7799, 7799, 
    7799, 7799, 7799, 8420, 8458, 8548, 8548, 8548, 8548, 8548,
  7700, 7851, 7761, 7775, 7786, 7793, 7801, 7806, 7812, 7829, 7829, 7829, 
    7829, 7829, 7829, 8411, 8459, 8547, 8547, 8547, 8547, 8547,
  7734, 7883, 7812, 7826, 7836, 7844, 7851, 7856, 7862, 7878, 7878, 7878, 
    7878, 7878, 7878, 8429, 8490, 8576, 8576, 8576, 8576, 8576,
  7773, 7931, 7968, 7982, 7993, 8001, 8009, 8013, 8020, 8036, 8036, 8036, 
    8036, 8036, 8036, 8484, 8625, 8708, 8708, 8708, 8708, 8708,
  7930, 8077, 8134, 8146, 8156, 8163, 8170, 8173, 8179, 8193, 8193, 8193, 
    8193, 8193, 8193, 8566, 8709, 8786, 8786, 8786, 8786, 8786,
  8087, 8316, 8371, 8372, 8372, 8372, 8372, 8371, 8371, 8371, 8371, 8371, 
    8371, 8371, 8371, 8550, 8369, 8369, 8369, 8369, 8369, 8369,
  8192, 8398, 8437, 8433, 8431, 8428, 8426, 8424, 8423, 8419, 8419, 8419, 
    8419, 8419, 8419, 8494, 8266, 8266, 8266, 8266, 8266, 8266,
  8361, 8528, 8523, 8512, 8504, 8498, 8492, 8488, 8483, 8471, 8471, 8471, 
    8471, 8471, 8471, 8389, 8047, 8047, 8047, 8047, 8047, 8047,
  8564, 8716, 8704, 8686, 8674, 8664, 8655, 8648, 8641, 8621, 8621, 8621, 
    8621, 8621, 8621, 8424, 7943, 7943, 7943, 7943, 7943, 7943,
  8572, 8705, 8646, 8630, 8618, 8609, 8600, 8594, 8588, 8569, 8569, 8569, 
    8569, 8569, 8569, 8377, 7939, 7939, 7939, 7939, 7939, 7939,
  8486, 8662, 8725, 8705, 8691, 8680, 8669, 8662, 8654, 8631, 8631, 8631, 
    8631, 8631, 8631, 8403, 7865, 7865, 7865, 7865, 7865, 7865,
  8341, 8582, 8778, 8757, 8742, 8731, 8719, 8711, 8704, 8680, 8680, 8680, 
    8680, 8680, 8680, 8501, 7873, 7873, 7873, 7873, 7873, 7873,
  8086, 8360, 8650, 8631, 8617, 8607, 8596, 8589, 8582, 8560, 8560, 8560, 
    8560, 8560, 8560, 8405, 7822, 7822, 7822, 7822, 7822, 7822,
  8838, 8940, 9058, 9050, 9045, 9042, 9039, 9036, 9034, 9026, 9026, 9026, 
    9026, 9026, 9026, 8963, 8772, 8772, 8772, 8772, 8772, 8772,
  8870, 8968, 8991, 8985, 8981, 8977, 8975, 8973, 8971, 8964, 8964, 8964, 
    8964, 8964, 8964, 8939, 8749, 8749, 8749, 8749, 8749, 8749,
  9026, 9117, 8970, 8967, 8964, 8962, 8962, 8960, 8959, 8955, 8955, 8955, 
    8955, 8955, 8955, 9003, 8834, 8834, 8834, 8834, 8834, 8834,
  8870, 8968, 8845, 8842, 8840, 8839, 8839, 8838, 8837, 8834, 8834, 8834, 
    8834, 8834, 8834, 8905, 8750, 8750, 8750, 8750, 8750, 8750,
  8533, 8657, 8580, 8582, 8583, 8585, 8587, 8587, 8588, 8591, 8591, 8591, 
    8591, 8591, 8591, 8771, 8682, 8682, 8682, 8682, 8682, 8682,
  9061, 9147, 9013, 9008, 9005, 9002, 9000, 8998, 8997, 8991, 8991, 8991, 
    8991, 8991, 8991, 9004, 8808, 8808, 8808, 8808, 8808, 8808,
  9157, 9235, 9200, 9186, 9176, 9169, 9163, 9158, 9153, 9138, 9138, 9138, 
    9138, 9138, 9138, 9020, 8635, 8635, 8635, 8635, 8635, 8635,
  8958, 9054, 8980, 8976, 8973, 8971, 8970, 8968, 8967, 8962, 8962, 8962, 
    8962, 8962, 8962, 8993, 8819, 8819, 8819, 8819, 8819, 8819,
  8903, 9005, 8941, 8936, 8932, 8930, 8928, 8927, 8925, 8919, 8919, 8919, 
    8919, 8919, 8919, 8963, 8751, 8751, 8751, 8751, 8751, 8751,
  8912, 9016, 8890, 8886, 8883, 8881, 8880, 8879, 8878, 8874, 8874, 8874, 
    8874, 8874, 8874, 8965, 8746, 8746, 8746, 8746, 8746, 8746,
  8914, 9016, 8848, 8846, 8845, 8844, 8844, 8844, 8843, 8841, 8841, 8841, 
    8841, 8841, 8841, 8959, 8788, 8788, 8788, 8788, 8788, 8788,
  8928, 9028, 8841, 8839, 8838, 8837, 8837, 8836, 8835, 8833, 8833, 8833, 
    8833, 8833, 8833, 8953, 8771, 8771, 8771, 8771, 8771, 8771,
  8936, 9036, 8878, 8874, 8872, 8870, 8869, 8868, 8866, 8862, 8862, 8862, 
    8862, 8862, 8862, 8957, 8738, 8737, 8737, 8737, 8737, 8737,
  8992, 9097, 8954, 8953, 8953, 8952, 8953, 8953, 8952, 8952, 8952, 8952, 
    8952, 8952, 8952, 9080, 8935, 8935, 8935, 8935, 8935, 8935,
  8968, 9074, 8871, 8873, 8874, 8875, 8877, 8878, 8879, 8881, 8881, 8881, 
    8881, 8881, 8881, 9062, 8962, 8962, 8962, 8962, 8962, 8962,
  9038, 9137, 8905, 8901, 8899, 8897, 8896, 8895, 8894, 8890, 8890, 8890, 
    8890, 8890, 8890, 9017, 8766, 8766, 8766, 8766, 8766, 8766,
  9104, 9194, 8959, 8953, 8949, 8946, 8943, 8941, 8939, 8932, 8932, 8932, 
    8932, 8932, 8932, 9013, 8714, 8714, 8714, 8714, 8714, 8714,
  9112, 9205, 8953, 8948, 8945, 8943, 8941, 8939, 8938, 8932, 8932, 8932, 
    8932, 8932, 8932, 9044, 8764, 8764, 8764, 8764, 8764, 8764,
  9163, 9249, 8898, 8892, 8888, 8885, 8883, 8881, 8879, 8872, 8872, 8872, 
    8872, 8872, 8872, 8997, 8666, 8666, 8666, 8666, 8666, 8666,
  9153, 9236, 8870, 8864, 8860, 8856, 8854, 8852, 8850, 8844, 8844, 8844, 
    8844, 8844, 8844, 8962, 8633, 8633, 8633, 8633, 8633, 8633,
  9044, 9133, 8749, 8746, 8744, 8743, 8743, 8742, 8741, 8738, 8738, 8738, 
    8738, 8738, 8738, 8912, 8652, 8652, 8652, 8652, 8652, 8652,
  9081, 9171, 8831, 8826, 8823, 8821, 8820, 8818, 8816, 8812, 8812, 8812, 
    8812, 8812, 8812, 8952, 8659, 8659, 8659, 8659, 8659, 8659,
  9005, 9106, 8679, 8678, 8677, 8677, 8677, 8677, 8676, 8675, 8675, 8675, 
    8675, 8675, 8675, 8927, 8641, 8641, 8641, 8641, 8641, 8641,
  8959, 9066, 8685, 8688, 8690, 8692, 8695, 8696, 8697, 8701, 8701, 8701, 
    8701, 8701, 8701, 8984, 8837, 8837, 8837, 8837, 8837, 8837,
  9059, 9151, 8799, 8795, 8792, 8790, 8789, 8787, 8786, 8781, 8781, 8781, 
    8781, 8781, 8781, 8943, 8644, 8644, 8644, 8644, 8644, 8644,
  9123, 9214, 8922, 8917, 8914, 8911, 8910, 8908, 8906, 8901, 8901, 8901, 
    8901, 8901, 8901, 9026, 8731, 8731, 8731, 8731, 8731, 8731,
  9014, 9119, 8808, 8812, 8815, 8817, 8820, 8821, 8822, 8826, 8826, 8826, 
    8826, 8826, 8826, 9072, 8979, 8979, 8979, 8979, 8979, 8979,
  9033, 9138, 8756, 8758, 8760, 8761, 8764, 8764, 8765, 8768, 8768, 8768, 
    8768, 8768, 8768, 9038, 8873, 8873, 8873, 8873, 8873, 8873,
  8916, 9026, 8607, 8611, 8613, 8615, 8618, 8620, 8621, 8625, 8625, 8625, 
    8625, 8625, 8625, 8942, 8774, 8774, 8774, 8774, 8774, 8774,
  8906, 9017, 8594, 8599, 8603, 8606, 8609, 8611, 8613, 8618, 8618, 8618, 
    8618, 8618, 8618, 8947, 8814, 8814, 8814, 8814, 8814, 8814,
  8843, 8956, 8502, 8505, 8508, 8509, 8512, 8513, 8515, 8518, 8518, 8518, 
    8518, 8518, 8518, 8862, 8657, 8657, 8657, 8657, 8657, 8657,
  8786, 8903, 8497, 8502, 8505, 8507, 8510, 8512, 8514, 8519, 8519, 8519, 
    8519, 8519, 8519, 8857, 8695, 8695, 8695, 8695, 8695, 8695,
  8953, 9064, 8668, 8673, 8677, 8679, 8683, 8685, 8687, 8692, 8692, 8692, 
    8692, 8692, 8692, 9011, 8893, 8893, 8893, 8893, 8893, 8893,
  8921, 9026, 8687, 8688, 8689, 8690, 8691, 8692, 8692, 8694, 8694, 8694, 
    8694, 8694, 8694, 8932, 8753, 8753, 8753, 8753, 8753, 8753,
  9126, 9220, 9021, 9020, 9019, 9018, 9018, 9018, 9017, 9016, 9016, 9016, 
    9016, 9016, 9016, 9126, 8973, 8973, 8973, 8973, 8973, 8973,
  9311, 9391, 9093, 9086, 9081, 9078, 9075, 9072, 9070, 9062, 9062, 9062, 
    9062, 9062, 9062, 9130, 8810, 8810, 8810, 8810, 8810, 8810,
  9322, 9401, 8985, 8981, 8978, 8976, 8975, 8974, 8972, 8967, 8967, 8967, 
    8967, 8967, 8967, 9109, 8822, 8822, 8822, 8822, 8822, 8822,
  9543, 9612, 9255, 9246, 9240, 9235, 9231, 9228, 9225, 9215, 9215, 9215, 
    9215, 9215, 9215, 9262, 8888, 8888, 8888, 8888, 8888, 8888,
  9444, 9519, 9178, 9175, 9173, 9171, 9170, 9169, 9168, 9165, 9165, 9165, 
    9165, 9165, 9165, 9263, 9058, 9058, 9058, 9058, 9058, 9058,
  9339, 9421, 9162, 9159, 9158, 9156, 9156, 9155, 9154, 9151, 9151, 9151, 
    9151, 9151, 9151, 9237, 9068, 9068, 9068, 9068, 9068, 9068,
  9189, 9276, 9105, 9101, 9099, 9097, 9095, 9094, 9093, 9088, 9088, 9088, 
    9088, 9088, 9088, 9140, 8949, 8949, 8949, 8949, 8949, 8949,
  8984, 9080, 8792, 8787, 8784, 8781, 8780, 8778, 8776, 8770, 8770, 8770, 
    8770, 8770, 8770, 8906, 8595, 8595, 8595, 8595, 8595, 8595,
  8514, 8637, 8278, 8280, 8282, 8283, 8285, 8286, 8287, 8290, 8290, 8290, 
    8290, 8290, 8290, 8609, 8389, 8389, 8389, 8389, 8389, 8389,
  8583, 8706, 8436, 8434, 8433, 8432, 8432, 8431, 8430, 8428, 8428, 8428, 
    8428, 8428, 8428, 8678, 8368, 8368, 8368, 8368, 8368, 8368,
  8344, 8483, 8115, 8119, 8121, 8123, 8126, 8128, 8129, 8133, 8133, 8133, 
    8133, 8133, 8133, 8533, 8289, 8289, 8289, 8289, 8289, 8289,
  8035, 8197, 7860, 7874, 7884, 7891, 7900, 7904, 7909, 7925, 7925, 7925, 
    7925, 7925, 7925, 8464, 8462, 8462, 8462, 8462, 8461, 8462,
  7908, 8079, 7752, 7775, 7792, 7804, 7817, 7825, 7833, 7859, 7859, 7859, 
    7859, 7859, 7859, 8481, 8730, 8730, 8730, 8730, 8730, 8730,
  7849, 8020, 7656, 7683, 7702, 7717, 7732, 7742, 7752, 7782, 7782, 7782, 
    7782, 7782, 7782, 8447, 8817, 8817, 8817, 8817, 8817, 8817,
  7892, 8064, 7645, 7673, 7693, 7708, 7723, 7733, 7743, 7774, 7774, 7774, 
    7774, 7774, 7774, 8474, 8827, 8827, 8827, 8827, 8826, 8827,
  7951, 8120, 7753, 7782, 7802, 7817, 7834, 7844, 7854, 7886, 7886, 7886, 
    7886, 7886, 7886, 8555, 8978, 8978, 8978, 8978, 8978, 8978,
  7999, 8162, 7797, 7815, 7828, 7838, 7848, 7855, 7861, 7881, 7881, 7881, 
    7881, 7881, 7881, 8460, 8574, 8574, 8574, 8574, 8574, 8574,
  7918, 8090, 7746, 7774, 7793, 7807, 7823, 7832, 7842, 7872, 7872, 7872, 
    7872, 7872, 7872, 8530, 8903, 8903, 8903, 8903, 8903, 8903,
  7861, 8040, 7627, 7653, 7672, 7686, 7700, 7710, 7719, 7748, 7748, 7748, 
    7748, 7748, 7748, 8465, 8742, 8742, 8742, 8742, 8742, 8742,
  7561, 7727, 7589, 7606, 7618, 7627, 7636, 7641, 7649, 7668, 7668, 7668, 
    7668, 7668, 7668, 8370, 8392, 8488, 8488, 8488, 8488, 8488,
  7687, 7880, 7248, 7272, 7289, 7301, 7315, 7324, 7332, 7358, 7358, 7358, 
    7358, 7358, 7358, 8229, 8258, 8258, 8258, 8258, 8258, 8258,
  7292, 7463, 7316, 7335, 7348, 7358, 7368, 7374, 7382, 7403, 7403, 7403, 
    7403, 7403, 7403, 8165, 8213, 8316, 8316, 8316, 8316, 8316,
  7070, 7260, 7205, 7226, 7241, 7252, 7263, 7270, 7279, 7302, 7302, 7302, 
    7302, 7302, 7302, 8045, 8181, 8287, 8287, 8287, 8287, 8287,
  7002, 7207, 7124, 7146, 7163, 7175, 7187, 7195, 7204, 7230, 7230, 7230, 
    7230, 7230, 7230, 8059, 8174, 8284, 8284, 8284, 8284, 8284,
  7013, 7212, 7165, 7187, 7203, 7215, 7227, 7234, 7243, 7269, 7269, 7269, 
    7269, 7269, 7269, 8039, 8187, 8295, 8295, 8295, 8295, 8295,
  7067, 7279, 7382, 7404, 7421, 7433, 7445, 7452, 7461, 7487, 7487, 7487, 
    7487, 7487, 7487, 8113, 8364, 8466, 8466, 8466, 8466, 8466,
  7113, 7316, 7424, 7445, 7461, 7473, 7484, 7491, 7500, 7524, 7524, 7524, 
    7524, 7524, 7524, 8113, 8370, 8470, 8470, 8470, 8470, 8470,
  7241, 7428, 7497, 7516, 7530, 7541, 7551, 7557, 7565, 7588, 7588, 7588, 
    7588, 7588, 7588, 8158, 8374, 8471, 8471, 8471, 8471, 8471,
  7436, 7597, 7531, 7548, 7560, 7569, 7578, 7583, 7590, 7609, 7609, 7609, 
    7609, 7609, 7609, 8232, 8328, 8423, 8423, 8423, 8423, 8423,
  7586, 7740, 7644, 7659, 7671, 7679, 7687, 7692, 7699, 7716, 7716, 7716, 
    7716, 7716, 7716, 8331, 8395, 8488, 8488, 8488, 8488, 8488,
  7685, 7824, 7719, 7733, 7743, 7750, 7757, 7762, 7768, 7783, 7783, 7783, 
    7783, 7783, 7783, 8355, 8405, 8495, 8495, 8495, 8495, 8495,
  7765, 7895, 7761, 7773, 7782, 7789, 7796, 7800, 7805, 7820, 7820, 7820, 
    7820, 7820, 7820, 8385, 8409, 8497, 8497, 8497, 8497, 8497,
  7810, 7935, 7795, 7807, 7815, 7822, 7828, 7832, 7837, 7851, 7851, 7851, 
    7851, 7851, 7851, 8404, 8420, 8508, 8508, 8508, 8508, 8508,
  7759, 7896, 7679, 7692, 7702, 7710, 7717, 7721, 7727, 7743, 7743, 7743, 
    7743, 7743, 7743, 8427, 8380, 8473, 8473, 8473, 8473, 8473,
  7694, 7867, 7805, 7821, 7834, 7842, 7851, 7856, 7864, 7882, 7882, 7882, 
    7882, 7882, 7882, 8497, 8557, 8646, 8646, 8646, 8646, 8646,
  7518, 7705, 7746, 7764, 7778, 7787, 7797, 7803, 7811, 7831, 7831, 7831, 
    7831, 7831, 7831, 8393, 8552, 8643, 8643, 8643, 8643, 8643,
  7343, 7540, 7597, 7617, 7631, 7642, 7652, 7659, 7667, 7690, 7690, 7690, 
    7690, 7690, 7690, 8287, 8473, 8568, 8568, 8568, 8568, 8568,
  7117, 7317, 7288, 7310, 7326, 7337, 7348, 7355, 7364, 7389, 7389, 7389, 
    7389, 7389, 7389, 8119, 8263, 8367, 8367, 8367, 8367, 8367,
  6945, 7169, 7090, 7114, 7132, 7146, 7159, 7167, 7177, 7205, 7205, 7205, 
    7205, 7205, 7205, 8088, 8196, 8307, 8307, 8307, 8307, 8307,
  6927, 7138, 7055, 7078, 7095, 7108, 7120, 7128, 7138, 7165, 7165, 7165, 
    7165, 7165, 7165, 8019, 8135, 8246, 8246, 8246, 8246, 8246,
  7050, 7254, 7091, 7114, 7130, 7142, 7154, 7162, 7171, 7197, 7197, 7197, 
    7197, 7197, 7197, 8104, 8143, 8253, 8253, 8253, 8253, 8253,
  7238, 7443, 7334, 7356, 7371, 7383, 7394, 7402, 7411, 7435, 7435, 7435, 
    7435, 7435, 7435, 8256, 8314, 8418, 8418, 8418, 8418, 8418,
  7441, 7633, 7526, 7546, 7560, 7570, 7581, 7587, 7595, 7618, 7618, 7618, 
    7618, 7618, 7618, 8371, 8412, 8510, 8510, 8510, 8510, 8510,
  7584, 7764, 7656, 7674, 7687, 7697, 7706, 7712, 7719, 7740, 7740, 7740, 
    7740, 7740, 7740, 8441, 8470, 8564, 8564, 8564, 8564, 8564,
  7614, 7798, 7669, 7687, 7700, 7710, 7720, 7726, 7733, 7754, 7754, 7754, 
    7754, 7754, 7754, 8487, 8495, 8589, 8589, 8589, 8589, 8589,
  7689, 7865, 7672, 7689, 7701, 7711, 7720, 7725, 7733, 7752, 7752, 7752, 
    7752, 7752, 7752, 8522, 8473, 8567, 8567, 8567, 8567, 8567,
  7722, 7882, 7689, 7705, 7716, 7724, 7733, 7738, 7744, 7762, 7762, 7762, 
    7762, 7762, 7762, 8481, 8436, 8528, 8528, 8528, 8528, 8528,
  7722, 7884, 7746, 7761, 7773, 7781, 7789, 7794, 7801, 7819, 7819, 7819, 
    7819, 7819, 7819, 8484, 8482, 8572, 8572, 8572, 8572, 8572,
  7662, 7821, 7706, 7722, 7733, 7741, 7750, 7755, 7761, 7779, 7779, 7779, 
    7779, 7779, 7779, 8417, 8443, 8534, 8534, 8534, 8534, 8534,
  7717, 7886, 7807, 7823, 7835, 7843, 7852, 7857, 7864, 7882, 7882, 7882, 
    7882, 7882, 7882, 8499, 8543, 8632, 8632, 8632, 8632, 8632,
  7704, 7870, 7839, 7855, 7866, 7875, 7883, 7888, 7895, 7913, 7913, 7913, 
    7913, 7913, 7913, 8471, 8557, 8645, 8645, 8645, 8645, 8645,
  7698, 7874, 7834, 7850, 7863, 7872, 7881, 7886, 7893, 7912, 7912, 7912, 
    7912, 7912, 7912, 8512, 8585, 8674, 8674, 8674, 8674, 8674,
  7773, 7945, 7905, 7921, 7933, 7941, 7950, 7955, 7962, 7980, 7980, 7980, 
    7980, 7980, 7980, 8554, 8620, 8706, 8706, 8706, 8706, 8706,
  7922, 8085, 8145, 8159, 8170, 8177, 8185, 8189, 8196, 8211, 8211, 8211, 
    8211, 8211, 8211, 8626, 8761, 8840, 8840, 8840, 8840, 8840,
  8061, 8197, 8238, 8249, 8258, 8263, 8269, 8273, 8278, 8290, 8290, 8290, 
    8290, 8290, 8290, 8632, 8750, 8824, 8824, 8824, 8824, 8824,
  8200, 8417, 8488, 8483, 8479, 8476, 8473, 8471, 8469, 8463, 8463, 8463, 
    8463, 8463, 8463, 8524, 8257, 8256, 8256, 8256, 8257, 8257,
  8405, 8582, 8606, 8594, 8585, 8578, 8571, 8566, 8562, 8547, 8547, 8547, 
    8547, 8547, 8547, 8447, 8066, 8066, 8066, 8066, 8066, 8066,
  8636, 8772, 8731, 8713, 8700, 8691, 8681, 8674, 8667, 8647, 8647, 8647, 
    8647, 8647, 8647, 8426, 7956, 7956, 7956, 7956, 7956, 7956,
  8569, 8694, 8670, 8648, 8632, 8620, 8608, 8600, 8592, 8567, 8567, 8567, 
    8567, 8567, 8567, 8249, 7721, 7721, 7721, 7721, 7721, 7721,
  8654, 8823, 8920, 8890, 8870, 8854, 8839, 8828, 8817, 8784, 8784, 8784, 
    8784, 8784, 8784, 8397, 7679, 7679, 7679, 7679, 7679, 7679,
  8443, 8652, 8807, 8780, 8762, 8748, 8734, 8724, 8714, 8684, 8684, 8684, 
    8684, 8684, 8684, 8392, 7684, 7684, 7684, 7684, 7684, 7684,
  8292, 8559, 8843, 8816, 8798, 8784, 8771, 8761, 8751, 8722, 8722, 8722, 
    8722, 8722, 8722, 8476, 7740, 7740, 7740, 7740, 7740, 7740,
  8862, 8968, 9138, 9130, 9125, 9121, 9119, 9116, 9114, 9106, 9106, 9106, 
    9106, 9106, 9106, 9035, 8850, 8850, 8850, 8850, 8850, 8850,
  8836, 8942, 8969, 8965, 8963, 8961, 8960, 8959, 8957, 8954, 8954, 8954, 
    8954, 8954, 8954, 8975, 8833, 8833, 8833, 8833, 8833, 8833,
  9141, 9237, 9228, 9214, 9204, 9196, 9189, 9184, 9179, 9163, 9163, 9163, 
    9163, 9163, 9163, 9103, 8634, 8634, 8634, 8634, 8634, 8634,
  8861, 8962, 8814, 8813, 8812, 8811, 8811, 8811, 8811, 8809, 8809, 8809, 
    8809, 8809, 8809, 8915, 8775, 8775, 8775, 8775, 8775, 8775,
  8966, 9058, 8941, 8936, 8933, 8931, 8929, 8928, 8926, 8921, 8921, 8921, 
    8921, 8921, 8921, 8955, 8756, 8756, 8756, 8756, 8756, 8756,
  9191, 9269, 9241, 9231, 9224, 9218, 9214, 9210, 9206, 9195, 9195, 9195, 
    9195, 9195, 9195, 9095, 8821, 8821, 8821, 8821, 8821, 8821,
  9026, 9121, 8986, 8985, 8984, 8984, 8984, 8984, 8984, 8983, 8983, 8983, 
    8983, 8983, 8983, 9064, 8958, 8958, 8958, 8958, 8958, 8958,
  8995, 9093, 8965, 8965, 8964, 8964, 8965, 8964, 8964, 8964, 8964, 8964, 
    8964, 8964, 8964, 9052, 8954, 8954, 8954, 8954, 8954, 8954,
  8886, 8988, 8910, 8906, 8904, 8902, 8901, 8899, 8898, 8893, 8893, 8893, 
    8893, 8893, 8893, 8954, 8758, 8758, 8758, 8758, 8758, 8758,
  9001, 9098, 8857, 8856, 8855, 8854, 8854, 8853, 8853, 8851, 8851, 8851, 
    8851, 8851, 8851, 8990, 8806, 8806, 8806, 8806, 8806, 8806,
  8920, 9020, 8853, 8851, 8850, 8849, 8849, 8849, 8848, 8846, 8846, 8846, 
    8846, 8846, 8846, 8956, 8788, 8788, 8788, 8788, 8788, 8788,
  8867, 8970, 8783, 8781, 8780, 8779, 8779, 8778, 8778, 8776, 8776, 8776, 
    8776, 8776, 8776, 8906, 8719, 8719, 8719, 8719, 8719, 8719,
  8979, 9083, 8971, 8970, 8970, 8969, 8970, 8969, 8969, 8968, 8968, 8968, 
    8968, 8968, 8968, 9075, 8947, 8947, 8947, 8947, 8947, 8947,
  8976, 9084, 8949, 8948, 8947, 8947, 8947, 8947, 8947, 8946, 8946, 8946, 
    8946, 8946, 8946, 9084, 8927, 8927, 8927, 8927, 8927, 8927,
  8939, 9048, 8876, 8874, 8873, 8872, 8873, 8872, 8872, 8870, 8870, 8870, 
    8870, 8870, 8870, 9024, 8826, 8826, 8826, 8826, 8826, 8826,
  9045, 9142, 8909, 8906, 8903, 8901, 8900, 8899, 8898, 8894, 8894, 8894, 
    8894, 8894, 8894, 9017, 8771, 8771, 8771, 8771, 8771, 8771,
  9118, 9206, 8972, 8966, 8962, 8959, 8956, 8954, 8952, 8946, 8946, 8946, 
    8946, 8946, 8946, 9018, 8736, 8736, 8736, 8736, 8736, 8736,
  9140, 9235, 9009, 9006, 9003, 9002, 9001, 9000, 8999, 8995, 8995, 8995, 
    8995, 8995, 8995, 9109, 8883, 8883, 8883, 8883, 8883, 8883,
  9154, 9246, 8988, 8984, 8982, 8980, 8979, 8978, 8976, 8972, 8972, 8972, 
    8972, 8972, 8972, 9089, 8852, 8852, 8852, 8852, 8852, 8852,
  9102, 9185, 8819, 8816, 8814, 8812, 8811, 8810, 8809, 8805, 8805, 8805, 
    8805, 8805, 8805, 8938, 8690, 8690, 8690, 8690, 8690, 8690,
  9051, 9141, 8774, 8771, 8769, 8768, 8767, 8766, 8765, 8762, 8762, 8762, 
    8762, 8762, 8762, 8923, 8661, 8661, 8661, 8661, 8661, 8661,
  9160, 9246, 8877, 8872, 8869, 8866, 8864, 8863, 8861, 8856, 8856, 8856, 
    8856, 8856, 8856, 8997, 8685, 8685, 8685, 8685, 8685, 8685,
  9099, 9195, 8748, 8745, 8743, 8742, 8742, 8741, 8740, 8737, 8737, 8737, 
    8737, 8737, 8737, 8973, 8650, 8650, 8650, 8650, 8650, 8650,
  9246, 9333, 8914, 8911, 8908, 8906, 8905, 8903, 8902, 8898, 8898, 8898, 
    8898, 8898, 8898, 9076, 8763, 8763, 8764, 8764, 8763, 8763,
  9156, 9244, 8889, 8884, 8881, 8878, 8876, 8875, 8873, 8867, 8867, 8867, 
    8867, 8867, 8867, 9004, 8691, 8691, 8691, 8691, 8691, 8691,
  9151, 9246, 8914, 8914, 8914, 8914, 8916, 8916, 8916, 8916, 8916, 8916, 
    8916, 8916, 8916, 9109, 8936, 8936, 8936, 8936, 8936, 8936,
  9157, 9250, 8884, 8885, 8885, 8886, 8887, 8888, 8888, 8889, 8889, 8889, 
    8889, 8889, 8889, 9094, 8934, 8934, 8934, 8934, 8934, 8934,
  9186, 9269, 8803, 8800, 8798, 8796, 8795, 8794, 8793, 8789, 8789, 8789, 
    8789, 8789, 8789, 8974, 8672, 8672, 8672, 8672, 8672, 8672,
  9127, 9214, 8818, 8816, 8815, 8814, 8813, 8813, 8812, 8809, 8809, 8809, 
    8809, 8809, 8809, 8979, 8737, 8737, 8737, 8737, 8737, 8737,
  8837, 8939, 8676, 8675, 8674, 8674, 8674, 8674, 8673, 8672, 8672, 8672, 
    8672, 8672, 8672, 8844, 8644, 8644, 8644, 8644, 8644, 8644,
  8775, 8891, 8639, 8641, 8641, 8642, 8643, 8644, 8644, 8645, 8645, 8645, 
    8645, 8645, 8645, 8879, 8696, 8696, 8696, 8696, 8696, 8696,
  8847, 8958, 8641, 8642, 8642, 8643, 8645, 8645, 8645, 8646, 8646, 8646, 
    8646, 8646, 8646, 8899, 8697, 8697, 8697, 8697, 8697, 8697,
  8805, 8916, 8522, 8522, 8522, 8522, 8523, 8523, 8523, 8522, 8522, 8522, 
    8522, 8522, 8522, 8804, 8528, 8528, 8528, 8528, 8528, 8528,
  8853, 8961, 8549, 8548, 8547, 8546, 8546, 8546, 8545, 8543, 8543, 8543, 
    8543, 8543, 8543, 8814, 8494, 8494, 8494, 8494, 8494, 8494,
  8790, 8898, 8640, 8640, 8640, 8641, 8642, 8642, 8642, 8642, 8642, 8642, 
    8642, 8642, 8642, 8840, 8667, 8667, 8667, 8667, 8667, 8667,
  8968, 9064, 8800, 8798, 8797, 8796, 8797, 8796, 8795, 8794, 8794, 8794, 
    8794, 8794, 8794, 8937, 8746, 8746, 8746, 8746, 8746, 8746,
  9252, 9332, 8974, 8970, 8967, 8965, 8964, 8962, 8961, 8956, 8956, 8956, 
    8956, 8956, 8956, 9075, 8810, 8810, 8810, 8810, 8810, 8810,
  9425, 9497, 9132, 9128, 9125, 9123, 9121, 9120, 9118, 9113, 9113, 9113, 
    9113, 9113, 9113, 9203, 8961, 8961, 8961, 8961, 8961, 8961,
  9489, 9559, 9221, 9212, 9206, 9202, 9198, 9195, 9193, 9183, 9183, 9183, 
    9183, 9183, 9183, 9225, 8882, 8882, 8882, 8882, 8882, 8882,
  9151, 9241, 8873, 8871, 8869, 8868, 8868, 8867, 8866, 8864, 8864, 8864, 
    8864, 8864, 8864, 9036, 8794, 8794, 8794, 8794, 8794, 8794,
  8938, 9039, 8729, 8728, 8728, 8727, 8728, 8728, 8728, 8727, 8727, 8727, 
    8727, 8727, 8727, 8920, 8718, 8718, 8718, 8718, 8718, 8718,
  8841, 8945, 8656, 8655, 8655, 8655, 8656, 8656, 8655, 8655, 8655, 8655, 
    8655, 8655, 8655, 8851, 8654, 8654, 8654, 8654, 8654, 8654,
  8562, 8689, 8445, 8448, 8449, 8451, 8453, 8454, 8455, 8457, 8457, 8457, 
    8457, 8457, 8457, 8738, 8559, 8559, 8559, 8559, 8559, 8559,
  8283, 8424, 8069, 8073, 8076, 8078, 8081, 8082, 8084, 8088, 8088, 8088, 
    8088, 8088, 8088, 8486, 8248, 8248, 8248, 8248, 8248, 8248,
  7974, 8139, 7746, 7761, 7771, 7779, 7788, 7793, 7799, 7815, 7815, 7815, 
    7815, 7815, 7815, 8401, 8384, 8384, 8384, 8384, 8384, 8384,
  7696, 7874, 7560, 7586, 7605, 7619, 7634, 7643, 7652, 7682, 7682, 7682, 
    7682, 7682, 7682, 8337, 8678, 8678, 8678, 8678, 8678, 8678,
  7645, 7827, 7461, 7489, 7508, 7522, 7537, 7547, 7556, 7587, 7587, 7587, 
    7587, 7587, 7587, 8293, 8612, 8612, 8612, 8612, 8612, 8612,
  7813, 7987, 7616, 7638, 7653, 7665, 7677, 7685, 7693, 7717, 7717, 7717, 
    7717, 7717, 7717, 8361, 8544, 8544, 8544, 8544, 8544, 8544,
  7701, 7814, 7719, 7730, 7739, 7745, 7751, 7754, 7759, 7772, 7772, 7772, 
    7772, 7772, 7772, 8257, 8331, 8418, 8418, 8418, 8418, 8418,
  7824, 7924, 7849, 7858, 7865, 7870, 7875, 7878, 7882, 7893, 7893, 7893, 
    7893, 7893, 7893, 8300, 8382, 8464, 8464, 8464, 8464, 8464,
  8087, 8249, 7844, 7856, 7865, 7871, 7879, 7883, 7887, 7901, 7901, 7901, 
    7901, 7901, 7901, 8460, 8367, 8367, 8367, 8367, 8367, 8367,
  7766, 7885, 7786, 7797, 7805, 7811, 7817, 7821, 7826, 7839, 7839, 7839, 
    7839, 7839, 7839, 8331, 8389, 8475, 8475, 8475, 8475, 8475,
  7565, 7690, 7564, 7577, 7586, 7593, 7600, 7604, 7610, 7625, 7625, 7625, 
    7625, 7625, 7625, 8194, 8253, 8346, 8346, 8346, 8346, 8346,
  7310, 7447, 7301, 7316, 7327, 7336, 7344, 7349, 7355, 7373, 7373, 7373, 
    7373, 7373, 7373, 8036, 8105, 8206, 8206, 8206, 8206, 8206,
  7152, 7302, 7124, 7141, 7154, 7163, 7172, 7178, 7185, 7205, 7205, 7205, 
    7205, 7205, 7205, 7965, 8019, 8126, 8126, 8126, 8126, 8126,
  6977, 7149, 7016, 7035, 7050, 7061, 7071, 7078, 7086, 7109, 7109, 7109, 
    7109, 7109, 7109, 7904, 8006, 8117, 8117, 8117, 8117, 8117,
  6857, 7060, 7045, 7068, 7085, 7097, 7109, 7117, 7126, 7152, 7152, 7152, 
    7152, 7152, 7152, 7917, 8110, 8221, 8221, 8221, 8221, 8221,
  6837, 7041, 6987, 7010, 7027, 7039, 7052, 7059, 7069, 7096, 7096, 7096, 
    7096, 7096, 7096, 7910, 8072, 8186, 8186, 8186, 8186, 8186,
  6916, 7123, 7164, 7187, 7203, 7216, 7228, 7235, 7245, 7271, 7271, 7271, 
    7271, 7271, 7271, 7973, 8198, 8305, 8305, 8305, 8305, 8305,
  7029, 7238, 7355, 7377, 7394, 7406, 7417, 7425, 7434, 7459, 7459, 7459, 
    7459, 7459, 7459, 8067, 8338, 8441, 8441, 8441, 8441, 8441,
  7211, 7413, 7493, 7514, 7529, 7541, 7552, 7559, 7567, 7591, 7591, 7591, 
    7591, 7591, 7591, 8196, 8417, 8515, 8515, 8515, 8515, 8515,
  7401, 7573, 7577, 7594, 7607, 7617, 7626, 7632, 7639, 7659, 7659, 7659, 
    7659, 7659, 7659, 8237, 8388, 8483, 8483, 8483, 8483, 8483,
  7555, 7711, 7673, 7688, 7700, 7708, 7716, 7721, 7728, 7745, 7745, 7745, 
    7745, 7745, 7745, 8302, 8411, 8501, 8501, 8501, 8501, 8501,
  7684, 7827, 7731, 7744, 7755, 7762, 7770, 7774, 7780, 7796, 7796, 7796, 
    7796, 7796, 7796, 8369, 8427, 8517, 8517, 8517, 8517, 8517,
  7775, 7893, 7767, 7778, 7787, 7793, 7799, 7803, 7808, 7821, 7821, 7821, 
    7821, 7821, 7821, 8343, 8379, 8466, 8466, 8466, 8466, 8466,
  7836, 7940, 7721, 7731, 7738, 7744, 7749, 7752, 7757, 7768, 7768, 7768, 
    7768, 7768, 7768, 8346, 8309, 8397, 8397, 8397, 8397, 8397,
  7854, 7957, 7752, 7761, 7769, 7774, 7779, 7782, 7787, 7798, 7798, 7798, 
    7798, 7798, 7798, 8358, 8330, 8416, 8416, 8416, 8416, 8416,
  7777, 7902, 7698, 7710, 7720, 7726, 7733, 7736, 7742, 7756, 7756, 7756, 
    7756, 7756, 7756, 8388, 8357, 8448, 8448, 8448, 8448, 8448,
  7675, 7847, 7786, 7802, 7815, 7824, 7832, 7838, 7845, 7864, 7864, 7864, 
    7864, 7864, 7864, 8478, 8540, 8630, 8630, 8630, 8630, 8630,
  7425, 7604, 7655, 7673, 7686, 7696, 7705, 7711, 7718, 7739, 7739, 7739, 
    7739, 7739, 7739, 8279, 8461, 8553, 8553, 8553, 8553, 8553,
  7208, 7413, 7436, 7457, 7473, 7484, 7495, 7502, 7511, 7536, 7536, 7536, 
    7536, 7536, 7536, 8209, 8379, 8480, 8480, 8480, 8480, 8480,
  7038, 7249, 7134, 7158, 7174, 7187, 7199, 7207, 7216, 7242, 7242, 7242, 
    7242, 7242, 7242, 8111, 8188, 8298, 8298, 8298, 8298, 8298,
  6880, 7093, 6890, 6914, 6931, 6945, 6957, 6965, 6975, 7003, 7003, 7003, 
    7003, 7003, 7003, 8001, 8026, 8143, 8143, 8143, 8143, 8143,
  6934, 7152, 7006, 7030, 7048, 7061, 7074, 7082, 7092, 7120, 7120, 7120, 
    7120, 7120, 7120, 8061, 8122, 8236, 8236, 8236, 8236, 8236,
  7105, 7326, 7204, 7227, 7245, 7258, 7270, 7278, 7288, 7315, 7315, 7315, 
    7315, 7315, 7315, 8214, 8269, 8378, 8378, 8378, 8378, 8378,
  7300, 7499, 7430, 7450, 7465, 7477, 7487, 7494, 7503, 7526, 7526, 7526, 
    7526, 7526, 7526, 8276, 8363, 8464, 8464, 8464, 8464, 8464,
  7508, 7694, 7639, 7657, 7671, 7681, 7691, 7697, 7704, 7725, 7725, 7725, 
    7725, 7725, 7725, 8392, 8470, 8564, 8564, 8564, 8564, 8564,
  7630, 7817, 7764, 7782, 7795, 7805, 7815, 7820, 7828, 7849, 7849, 7849, 
    7849, 7849, 7849, 8502, 8566, 8657, 8657, 8657, 8657, 8657,
  7700, 7876, 7737, 7754, 7767, 7776, 7785, 7790, 7797, 7817, 7817, 7817, 
    7817, 7817, 7817, 8525, 8517, 8609, 8609, 8609, 8609, 8609,
  7781, 7938, 7765, 7780, 7791, 7799, 7807, 7812, 7818, 7835, 7835, 7835, 
    7835, 7835, 7835, 8517, 8484, 8574, 8574, 8574, 8574, 8574,
  7771, 7921, 7636, 7651, 7662, 7670, 7678, 7682, 7689, 7706, 7706, 7706, 
    7706, 7706, 7706, 8497, 8381, 8475, 8475, 8475, 8475, 8475,
  7731, 7899, 7778, 7794, 7806, 7814, 7823, 7828, 7835, 7853, 7853, 7853, 
    7853, 7853, 7853, 8513, 8522, 8612, 8612, 8612, 8612, 8612,
  7687, 7857, 7749, 7765, 7777, 7786, 7794, 7800, 7807, 7825, 7825, 7825, 
    7825, 7825, 7825, 8481, 8504, 8595, 8595, 8595, 8595, 8595,
  7687, 7868, 7803, 7821, 7833, 7843, 7852, 7857, 7865, 7884, 7884, 7884, 
    7884, 7884, 7884, 8523, 8574, 8664, 8664, 8664, 8664, 8664,
  7710, 7888, 7883, 7900, 7912, 7921, 7930, 7935, 7943, 7961, 7961, 7961, 
    7961, 7961, 7961, 8522, 8621, 8708, 8708, 8708, 8708, 8708,
  7696, 7877, 7889, 7906, 7918, 7927, 7936, 7942, 7949, 7968, 7968, 7968, 
    7968, 7968, 7968, 8518, 8632, 8719, 8719, 8719, 8719, 8719,
  7735, 7906, 7915, 7931, 7943, 7952, 7960, 7965, 7972, 7990, 7990, 7990, 
    7990, 7990, 7990, 8514, 8625, 8711, 8711, 8711, 8711, 8711,
  7890, 8056, 8146, 8160, 8171, 8179, 8187, 8191, 8198, 8214, 8214, 8214, 
    8214, 8214, 8214, 8606, 8770, 8848, 8848, 8848, 8848, 8848,
  8038, 8195, 8277, 8290, 8299, 8306, 8313, 8317, 8323, 8338, 8338, 8338, 
    8338, 8338, 8338, 8696, 8838, 8912, 8912, 8912, 8912, 8912,
  8187, 8410, 8492, 8489, 8487, 8485, 8483, 8481, 8480, 8476, 8476, 8476, 
    8476, 8476, 8476, 8564, 8339, 8339, 8339, 8339, 8339, 8339,
  8463, 8662, 8709, 8695, 8685, 8677, 8670, 8664, 8659, 8643, 8643, 8643, 
    8643, 8643, 8643, 8574, 8101, 8101, 8101, 8101, 8101, 8102,
  8681, 8858, 8892, 8871, 8857, 8847, 8836, 8829, 8821, 8799, 8799, 8799, 
    8799, 8799, 8799, 8606, 8039, 8039, 8039, 8039, 8039, 8039,
  8699, 8838, 8796, 8776, 8762, 8751, 8741, 8733, 8726, 8704, 8704, 8704, 
    8704, 8704, 8704, 8478, 7953, 7953, 7953, 7953, 7953, 7953,
  8717, 8863, 8906, 8878, 8859, 8844, 8829, 8819, 8809, 8778, 8778, 8778, 
    8778, 8778, 8778, 8393, 7732, 7732, 7732, 7732, 7732, 7732,
  8548, 8757, 8934, 8904, 8884, 8868, 8852, 8842, 8831, 8798, 8798, 8798, 
    8798, 8798, 8798, 8444, 7684, 7684, 7684, 7684, 7684, 7684,
  8325, 8561, 8815, 8786, 8766, 8750, 8735, 8724, 8714, 8681, 8681, 8681, 
    8681, 8681, 8681, 8335, 7584, 7584, 7584, 7584, 7584, 7585 ;

 Freq = 23.8, 31.4, 50.3, 51.76, 52.8, 53.596, 54.4, 54.94, 55.5, 57.29, 
    57.29, 57.29, 57.29, 57.29, 57.29, 88.2, 165.5, 183.31, 183.31, 183.31, 
    183.31, 183.31 ;

 GWP =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 22, 26, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 0, 0, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 25, 35, 18, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 6, 23, 17, 20, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 7, 33, 14, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 12, 26, 10, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, 0, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 5, 15, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 10, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 6, 13, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 8, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, _, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 6, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, 
    _, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 IWP =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 LWP =
  0, 0, 0, 0, 0, 0, 0, 0, 1, 25, 9, 13, 7, 9, 49, 36, 39, 20, 2, 3, 23, 30, 
    30, 39, 40, 34, 31, 29, 33, 39, 44, 40, 45, 61, 59, 52, 41, 32, 40, 36, 
    34, 19, 7, 10, 13, 8, 1, 8, 15, 7, 1, 4, 4, 4, 5, 5, 5, 7, 5, -998, -998, 
    -998, -998, -998, -998, -998, -998, -998, -998, -998, -998, -998, -998, 
    -998, -998, -998, -998, -998, -998, -998, -998, -998, -998, -998, -998, 
    -998, -998, -998, -998, 5, 5, -998, -998, -998, -998, -998,
  0, 0, 0, 0, 0, 0, 0, 2, 14, 9, 10, 10, 11, 8, 53, 51, 31, 31, 27, 34, 33, 
    47, 52, 57, 38, 40, 33, 39, 33, 38, 37, 38, 36, 37, 34, 50, 49, 59, 47, 
    36, 27, 23, 8, 6, 6, 7, 10, 7, 3, 1, 2, 2, 3, 3, 5, 3, 3, 5, 11, 9, -998, 
    -998, -998, -998, -998, -998, -998, -998, -998, -998, -998, -998, -998, 
    -998, -998, -998, -998, -998, -998, -998, -998, -998, -998, -998, -998, 
    -998, -998, -998, -998, -998, -998, -998, -998, -998, -998, -998,
  0, 0, 0, 0, 0, 0, 1, 23, 8, 14, 17, 13, 9, 54, 36, 66, 41, 32, 37, 28, 32, 
    33, 33, 32, 41, 51, 39, 38, 31, 9, 11, 17, 29, 36, 35, 34, 43, 36, 43, 
    39, 26, 24, 19, 9, 7, 6, 9, 10, 5, 1, 3, 3, 3, 4, 6, 3, 1, 3, 13, 13, 6, 
    -998, -998, -998, -998, -998, -998, -998, -998, -998, -998, -998, -998, 
    -998, -998, -998, -998, -998, -998, -998, -998, -998, -998, -998, -998, 
    -998, -998, -998, -998, -998, -998, -998, -998, -998, -998, -998,
  0, 0, 0, 0, 0, 1, 13, 36, 13, 10, 12, 11, 39, 37, 34, 38, 40, 44, 42, 33, 
    32, 44, 37, 44, 44, 38, 30, 48, 12, 25, 30, 36, 24, 39, 42, 39, 28, 28, 
    31, 33, 29, 26, 10, 7, 6, 9, 15, 21, 11, 5, 3, 2, 8, 5, 4, 4, 2, 2, 9, 
    12, 8, -998, -998, -998, -998, -998, -998, -998, -998, -998, -998, -998, 
    -998, -998, -998, -998, -998, -998, -998, -998, -998, -998, -998, -998, 
    -998, -998, -998, -998, -998, -998, -998, -998, -998, -998, -998, -998,
  0, 0, 0, 0, 0, 5, 17, 22, 15, 13, 13, 9, 54, 24, 26, 44, 41, 40, 34, 34, 
    37, 58, 109, 56, 37, 53, 45, 39, 12, 10, 8, 7, 12, 33, 16, 26, 14, 11, 
    24, 26, 25, 6, 3, 3, 4, 14, 32, 10, 8, 9, 15, 13, 5, 5, 5, 2, 5, 4, 5, 9, 
    9, -998, 0, -998, -998, -998, -998, -998, -998, -998, -998, -998, -998, 
    -998, -998, -998, -998, -998, -998, -998, -998, -998, -998, -998, -998, 
    -998, -998, -998, -998, -998, -998, -998, -998, -998, -998, -998,
  0, 3, 5, 1, 12, 1, 13, 10, 17, 13, 41, 107, 61, 41, 31, 32, 38, 33, 28, 31, 
    34, 59, 89, 35, 25, 36, 35, 40, 10, 7, 8, 6, 11, 13, 14, 28, 28, 10, 21, 
    26, 25, 6, 3, 4, 17, 7, 8, 6, 22, 33, 32, 8, 6, 3, 2, 6, 7, 7, 6, 11, 
    -998, -998, -998, -998, -998, -998, -998, -998, -998, -998, -998, -998, 
    -998, -998, -998, -998, -998, -998, -998, -998, -998, -998, -998, -998, 
    -998, -998, -998, -998, -998, -998, -998, -998, -998, -998, -998, -998,
  9, 19, 17, 17, 19, 11, 44, 12, 12, 38, 29, 67, 57, 30, 28, 35, 42, 30, 30, 
    66, 86, 71, 32, 45, 38, 31, 15, 24, 5, 4, 7, 8, 31, 38, 39, 33, 23, 11, 
    29, 28, 26, 15, 45, 71, 56, 55, 41, 23, 11, 8, 9, 5, 3, 1, 6, 4, 7, 10, 
    15, 8, -998, -998, -998, -998, -998, -998, -998, -998, -998, -998, -998, 
    -998, -998, -998, -998, -998, -998, -998, -998, -998, -998, -998, -998, 
    -998, -998, -998, -998, -998, -998, -998, -998, -998, -998, -998, -998, 
    -998,
  7, 15, 23, 23, 13, 51, 11, 11, 10, 32, 40, 37, 28, 4, 20, 25, 6, 25, 32, 
    65, 55, 41, 33, 35, 33, 8, 33, 29, 6, 7, 9, 8, 20, 38, 36, 32, 35, 24, 
    22, 28, 26, 77, 88, 82, 66, 53, 53, 29, 5, 5, 7, 3, 3, 2, 5, 7, 12, 17, 
    11, 1, -998, -998, -998, -998, -998, -998, -998, -998, -998, -998, -998, 
    -998, -998, -998, -998, -998, -998, -998, -998, -998, -998, -998, -998, 
    -998, -998, -998, -998, -998, -998, -998, -998, -998, -998, -998, -998, 
    -998,
  14, 5, 15, 22, 33, 10, 10, 65, 28, 10, 19, 24, 30, 6, 3, 8, 37, 32, 40, 
    100, 45, 37, 30, 33, 39, 12, 87, 31, 4, 5, 8, 6, 20, 34, 43, 39, 93, 76, 
    32, 66, 90, 69, 29, 30, 30, 29, 12, 6, 4, 2, 4, 3, 7, 6, 6, 10, 14, -998, 
    -998, -998, -998, -998, -998, -998, -998, -998, -998, -998, -998, -998, 
    -998, -998, -998, -998, -998, -998, -998, -998, -998, -998, -998, -998, 
    -998, -998, -998, -998, -998, -998, -998, -998, -998, -998, -998, -998, 
    -998, -998,
  8, 3, 17, 31, 76, 10, 36, 9, 2, 3, 15, 29, 27, 4, 6, 11, 30, 11, 23, 30, 
    29, 13, 35, 32, 9, 26, 31, 4, 4, 5, 5, 11, 14, 11, 11, 21, 60, 31, 18, 
    32, 43, 7, 43, 34, 14, 9, 6, 3, 5, 5, 4, 8, 11, 10, 1, 11, 13, -998, 
    -998, -998, -998, -998, -998, -998, -998, -998, -998, -998, -998, -998, 
    -998, -998, -998, -998, -998, -998, -998, -998, -998, -998, -998, -998, 
    -998, -998, -998, -998, -998, -998, -998, -998, -998, -998, -998, -998, 
    -998, -998,
  7, 6, 17, 49, 86, 28, 5, 1, 21, 24, 26, 28, 31, 6, 7, 14, 29, 14, 30, 34, 
    32, 41, 26, 6, 37, 28, 7, 6, 8, 6, 13, 11, 7, 9, 13, 24, 32, 9, 6, 5, 7, 
    35, 26, 20, 6, 3, 1, 0, 0, 1, 5, 2, 1, -998, 3, -998, -998, -998, -998, 
    -998, -998, -998, -998, -998, -998, -998, -998, -998, -998, -998, -998, 
    -998, -998, -998, -998, -998, -998, -998, -998, -998, -998, -998, -998, 
    -998, -998, -998, -998, -998, -998, -998, -998, -998, -998, -998, -998, 
    -998,
  14, 3, 9, 35, 30, 10, 3, 3, 26, 27, 25, 28, 9, 6, 8, 25, 35, 19, 15, 35, 
    28, 40, 25, 36, 45, 11, 7, 30, 36, 31, 19, 12, 8, 24, 39, 42, 28, 7, 34, 
    41, 46, 37, 13, 8, 3, 2, 2, 0, -998, -998, 0, -998, -998, -998, -998, 
    -998, -998, -998, -998, -998, -998, -998, -998, -998, -998, -998, -998, 
    -998, -998, -998, -998, -998, -998, -998, -998, -998, -998, -998, -998, 
    -998, -998, -998, -998, -998, -998, -998, -998, -998, -998, -998, -998, 
    -998, -998, -998, -998, -998 ;

 LZ_angle =
  -63.96, -62.26001, -60.59999, -58.96998, -57.40001, -55.88, -54.39001, 
    -52.90001, -51.43, -49.97999, -48.57, -47.16999, -45.77, -44.37, 
    -42.98999, -41.64001, -40.29999, -38.95001, -37.59999, -36.27, -34.96, 
    -33.65001, -32.33001, -31.01, -29.71, -28.42999, -27.16, -25.85999, 
    -24.56, -23.28, -22.01, -20.75, -19.47, -18.19, -16.92999, -15.67, 
    -14.41, -13.14, -11.87, -10.61, -9.369999, -8.119999, -6.86, -5.580001, 
    -4.339999, -3.099999, -1.86, -0.5900001, 0.6800001, 1.93, 3.18, 4.43, 
    5.699999, 6.970001, 8.22, 9.460003, 10.72, 11.99, 13.26, 14.51, 15.76, 
    17.02, 18.31, 19.6, 20.87, 22.13, 23.4, 24.7, 25.99, 27.27, 28.54999, 
    29.85, 31.16, 32.46999, 33.77, 35.07, 36.40999, 37.76001, 39.10999, 
    40.44, 41.77, 43.14001, 44.53001, 45.93, 47.32, 48.71999, 50.15001, 
    51.60999, 53.08001, 54.56001, 56.06001, 57.60999, 59.2, 60.83, 62.46998, 
    64.16003,
  -63.96998, -62.23999, -60.58, -58.97999, -57.43001, -55.89001, -54.37, 
    -52.89001, -51.43, -50.01001, -48.57, -47.15001, -45.73999, -44.37, 
    -43.01001, -41.65001, -40.28001, -38.93, -37.59999, -36.29999, -34.96999, 
    -33.63, -32.31, -31.01, -29.73, -28.44, -27.14001, -25.84, -24.57001, 
    -23.3, -22.02, -20.73, -19.45999, -18.2, -16.95, -15.67, -14.39, -13.12, 
    -11.88, -10.64, -9.369999, -8.11, -6.839998, -5.599999, -4.36, -3.099999, 
    -1.83, -0.58, 0.67, 1.91, 3.18, 4.46, 5.699999, 6.949998, 8.199998, 
    9.460003, 10.74, 11.99, 13.24, 14.49, 15.77, 17.05, 18.32001, 19.57999, 
    20.85, 22.13, 23.42001, 24.69, 25.97, 27.26, 28.56, 29.88, 31.17, 
    32.45001, 33.76001, 35.09001, 36.43, 37.76001, 39.08001, 40.41999, 
    41.78999, 43.16999, 44.53001, 45.90999, 47.31, 48.72999, 50.16999, 
    51.60999, 53.05, 54.55, 56.09, 57.64001, 59.2, 60.8, 62.46, 64.18999,
  -63.93999, -62.22999, -60.59999, -58.98999, -57.41, -55.87, -54.37, 
    -52.90001, -51.43, -49.97999, -48.53999, -47.14001, -45.77, -44.39001, 
    -43, -41.62, -40.27, -38.95001, -37.62, -36.28001, -34.96, -33.64001, 
    -32.34001, -31.03001, -29.71999, -28.41, -27.14001, -25.85999, -24.57999, 
    -23.28, -22, -20.74, -19.48, -18.22, -16.92999, -15.65, -14.4, -13.15, 
    -11.89, -10.61, -9.36, -8.11, -6.86, -5.61, -4.339999, -3.080001, -1.84, 
    -0.6000001, 0.6599999, 1.93, 3.2, 4.440001, 5.68, 6.940001, 8.22, 
    9.479997, 10.73, 11.98, 13.24, 14.52, 15.78, 17.03, 18.29001, 19.57999, 
    20.87, 22.14001, 23.4, 24.67999, 25.98, 27.28, 28.58, 29.85, 31.14001, 
    32.45001, 33.78001, 35.09999, 36.40999, 37.73999, 39.09001, 40.45001, 
    41.79999, 43.15001, 44.52, 45.91999, 47.33001, 48.72999, 50.15001, 
    51.59001, 53.07, 54.58001, 56.09, 57.62, 59.18999, 60.81001, 62.48999, 
    64.18999,
  -63.96998, -62.26001, -60.59, -58.96998, -57.41, -55.90001, -54.40001, 
    -52.90001, -51.41999, -49.97999, -48.57, -47.16999, -45.76001, -44.35999, 
    -42.98999, -41.64001, -40.29999, -38.94, -37.59001, -36.28001, -34.96999, 
    -33.65999, -32.33001, -31.01, -29.71, -28.44, -27.15, -25.85, -24.55, 
    -23.28, -22.02, -20.75, -19.47, -18.19, -16.92999, -15.67, -14.4, -13.13, 
    -11.86, -10.62, -9.380001, -8.119999, -6.85, -5.580001, -4.339999, 
    -3.099999, -1.85, -0.58, 0.6800001, 1.93, 3.169999, 4.43, 5.699999, 
    6.970001, 8.210002, 9.460003, 10.72, 12, 13.26, 14.51, 15.76, 17.03, 
    18.32001, 19.6, 20.85999, 22.13, 23.4, 24.7, 25.99, 27.27, 28.54999, 
    29.85, 31.17, 32.46999, 33.77, 35.08001, 36.41999, 37.77, 39.10999, 
    40.43, 41.78001, 43.15001, 44.53999, 45.93, 47.31, 48.71001, 50.15999, 
    51.62, 53.08001, 54.55, 56.07, 57.63, 59.21998, 60.83, 62.46, 64.17001,
  -63.95, -62.21998, -60.56999, -58.97999, -57.42, -55.88, -54.35999, -52.88, 
    -51.43, -50, -48.56, -47.13, -45.73999, -44.37, -43.02, -41.64001, 
    -40.27, -38.91999, -37.60999, -36.29, -34.96999, -33.63, -32.32, -31.02, 
    -29.73, -28.42999, -27.13, -25.84, -24.57001, -23.3, -22.01, -20.72, 
    -19.45999, -18.20999, -16.95, -15.67, -14.38, -13.13, -11.88, -10.64, 
    -9.369999, -8.100001, -6.839998, -5.61, -4.349999, -3.09, -1.83, -0.58, 
    0.6599999, 1.92, 3.19, 4.46, 5.699999, 6.940001, 8.199998, 9.47, 10.74, 
    12, 13.24, 14.5, 15.77, 17.05, 18.31, 19.57999, 20.85, 22.14001, 
    23.42001, 24.7, 25.97, 27.27, 28.57001, 29.87, 31.16, 32.45001, 33.76001, 
    35.09999, 36.43, 37.76001, 39.08001, 40.43, 41.79999, 43.16999, 44.53001, 
    45.90999, 47.32, 48.75, 50.18, 51.60999, 53.06001, 54.56001, 56.09999, 
    57.65001, 59.2, 60.8, 62.46998, 64.19999,
  -63.93001, -62.22999, -60.59, -58.98999, -57.41, -55.87, -54.38, -52.90999, 
    -51.43, -49.97999, -48.53999, -47.15001, -45.77, -44.38, -42.98999, 
    -41.62, -40.28001, -38.95001, -37.60999, -36.27, -34.95001, -33.64001, 
    -32.34001, -31.03001, -29.71, -28.42, -27.14001, -25.85999, -24.57001, 
    -23.27, -22, -20.74, -19.48, -18.20999, -16.92, -15.66, -14.4, -13.15, 
    -11.88, -10.61, -9.350002, -8.11, -6.86, -5.589998, -4.330001, -3.080001, 
    -1.85, -0.6000001, 0.67, 1.94, 3.2, 4.43, 5.68, 6.949998, 8.229997, 
    9.479997, 10.72, 11.98, 13.25, 14.53, 15.78, 17.03, 18.3, 19.59, 20.88, 
    22.14001, 23.4, 24.69, 25.98, 27.28, 28.56, 29.85, 31.15, 32.46999, 
    33.79, 35.09999, 36.40999, 37.73999, 39.09999, 40.45001, 41.78999, 
    43.15001, 44.53001, 45.93, 47.34001, 48.72999, 50.14001, 51.59999, 
    53.08001, 54.58001, 56.08001, 57.62, 59.2, 60.81999, 62.48999, 64.18999,
  -63.96998, -62.25, -60.59, -58.96998, -57.41, -55.90001, -54.39001, 
    -52.90001, -51.43, -49.98999, -48.58001, -47.16999, -45.75, -44.34999, 
    -43, -41.64001, -40.28999, -38.93, -37.59001, -36.28001, -34.96999, 
    -33.65001, -32.32, -31.01, -29.71999, -28.44, -27.15, -25.84, -24.55, 
    -23.29001, -22.02, -20.75, -19.47, -18.19, -16.94, -15.68, -14.4, -13.12, 
    -11.86, -10.62, -9.380001, -8.119999, -6.839998, -5.580001, -4.339999, 
    -3.099999, -1.84, -0.58, 0.6800001, 1.92, 3.18, 4.440001, 5.71, 6.960001, 
    8.210002, 9.460003, 10.73, 12, 13.26, 14.5, 15.76, 17.04001, 18.32999, 
    19.6, 20.85999, 22.13, 23.41, 24.7, 25.98, 27.26, 28.54999, 29.85999, 
    31.17, 32.46999, 33.76001, 35.08001, 36.41999, 37.77, 39.09999, 40.43, 
    41.78001, 43.15001, 44.53999, 45.91999, 47.31, 48.71999, 50.16999, 51.62, 
    53.08001, 54.55, 56.07, 57.63, 59.21998, 60.81001, 62.46, 64.18002,
  -63.95, -62.21998, -60.56999, -58.98999, -57.43001, -55.88, -54.37, 
    -52.89001, -51.43999, -50, -48.56, -47.13, -45.75, -44.38, -43.01001, 
    -41.63, -40.27, -38.93, -37.62, -36.29999, -34.96, -33.63, -32.32, 
    -31.03001, -29.73, -28.42999, -27.13, -25.85, -24.57001, -23.29001, -22, 
    -20.72, -19.47, -18.22, -16.94, -15.66, -14.39, -13.14, -11.89, -10.63, 
    -9.36, -8.100001, -6.85, -5.61, -4.349999, -3.09, -1.83, -0.5900001, 
    0.6499999, 1.92, 3.19, 4.449999, 5.690001, 6.940001, 8.210002, 9.479997, 
    10.75, 11.99, 13.24, 14.5, 15.78, 17.05, 18.31, 19.57999, 20.85999, 
    22.14001, 23.42001, 24.67999, 25.96, 27.26, 28.58, 29.87, 31.15, 
    32.45001, 33.77, 35.09999, 36.43, 37.73999, 39.08001, 40.43, 41.79999, 
    43.16999, 44.52, 45.90999, 47.32, 48.73999, 50.15999, 51.59001, 53.06001, 
    54.57, 56.09999, 57.65001, 59.18999, 60.8, 62.46998, 64.19999,
  -63.93999, -62.22999, -60.59, -58.96998, -57.40001, -55.87, -54.38, 
    -52.90999, -51.43, -49.96999, -48.54999, -47.15999, -45.77, -44.38, 
    -42.98, -41.62, -40.28999, -38.95001, -37.60999, -36.27, -34.96, 
    -33.65001, -32.34001, -31.02, -29.71999, -28.42999, -27.15, -25.85999, 
    -24.57001, -23.28, -22.01, -20.75, -19.49, -18.20999, -16.92999, -15.66, 
    -14.41, -13.15, -11.88, -10.61, -9.36, -8.119999, -6.86, -5.589998, 
    -4.330001, -3.09, -1.86, -0.6000001, 0.6800001, 1.95, 3.19, 4.43, 
    5.690001, 6.949998, 8.22, 9.47, 10.72, 11.98, 13.26, 14.52, 15.77, 17.02, 
    18.3, 19.59, 20.87, 22.13, 23.4, 24.67999, 25.99, 27.28, 28.56, 29.85, 
    31.15, 32.46999, 33.78001, 35.08001, 36.40999, 37.75, 39.10999, 40.45001, 
    41.78999, 43.14001, 44.53001, 45.93, 47.33001, 48.72999, 50.14001, 
    51.59999, 53.08001, 54.57, 56.08001, 57.60999, 59.2, 60.81999, 62.47999, 
    64.18002,
  -63.96998, -62.25, -60.58, -58.97999, -57.42, -55.90001, -54.39001, 
    -52.89001, -51.43999, -50, -48.58001, -47.15999, -45.75, -44.35999, 
    -43.01001, -41.65001, -40.28001, -38.93, -37.59999, -36.29, -34.98, 
    -33.65001, -32.32, -31.02, -29.73, -28.45001, -27.14001, -25.84, -24.56, 
    -23.29001, -22.02, -20.74, -19.45999, -18.20999, -16.95, -15.68, -14.4, 
    -13.13, -11.87, -10.63, -9.380001, -8.11, -6.839998, -5.589998, 
    -4.349999, -3.099999, -1.84, -0.58, 0.67, 1.92, 3.18, 4.449999, 5.71, 
    6.949998, 8.190001, 9.460003, 10.73, 12, 13.25, 14.49, 15.76, 17.04001, 
    18.32001, 19.59, 20.85, 22.13, 23.42001, 24.7, 25.98, 27.26, 28.56, 
    29.87, 31.17, 32.45001, 33.76001, 35.09001, 36.43, 37.77, 39.09001, 
    40.41999, 41.78001, 43.15999, 44.53999, 45.90999, 47.31, 48.72999, 
    50.16999, 51.62, 53.07, 54.55, 56.08001, 57.65001, 59.21, 60.8, 62.46, 
    64.18002,
  -63.93999, -62.21998, -60.58, -58.98999, -57.41, -55.87, -54.35999, 
    -52.89001, -51.43999, -49.98999, -48.54999, -47.14001, -45.76001, -44.38, 
    -43, -41.62, -40.26001, -38.94, -37.63, -36.29, -34.96, -33.63, 
    -32.33001, -31.03001, -29.73, -28.42, -27.13, -25.85999, -24.57999, 
    -23.29001, -22, -20.73, -19.47, -18.22, -16.94, -15.65, -14.39, -13.14, 
    -11.89, -10.63, -9.36, -8.100001, -6.86, -5.61, -4.349999, -3.080001, 
    -1.83, -0.6000001, 0.6599999, 1.93, 3.19, 4.449999, 5.690001, 6.940001, 
    8.210002, 9.479997, 10.73, 11.98, 13.24, 14.51, 15.78, 17.04001, 18.3, 
    19.57999, 20.85999, 22.14001, 23.42001, 24.67999, 25.97, 27.28, 28.58, 
    29.85999, 31.15, 32.45001, 33.77, 35.09999, 36.41999, 37.73999, 39.08001, 
    40.44, 41.79999, 43.15001, 44.52, 45.90999, 47.33001, 48.73999, 50.15999, 
    51.58001, 53.06001, 54.57, 56.09999, 57.63, 59.18999, 60.81001, 62.48999, 
    64.19999,
  -63.96, -62.26001, -60.60999, -58.97999, -57.41, -55.88, -54.39001, 
    -52.90999, -51.43, -49.97999, -48.56, -47.16999, -45.77, -44.37, 
    -42.98999, -41.64001, -40.28999, -38.95001, -37.59999, -36.27, -34.96, 
    -33.65001, -32.34001, -31.01, -29.71, -28.42999, -27.16, -25.85999, 
    -24.56, -23.28, -22.01, -20.75, -19.47, -18.2, -16.92999, -15.67, -14.41, 
    -13.14, -11.87, -10.62, -9.369999, -8.119999, -6.86, -5.580001, 
    -4.330001, -3.099999, -1.85, -0.6000001, 0.6800001, 1.94, 3.19, 4.43, 
    5.699999, 6.960001, 8.210002, 9.460003, 10.72, 11.99, 13.27, 14.52, 
    15.76, 17.02, 18.31, 19.6, 20.87, 22.12, 23.4, 24.7, 26, 27.28, 28.54999, 
    29.85, 31.16, 32.46999, 33.77, 35.08001, 36.40999, 37.76001, 39.10999, 
    40.44, 41.78001, 43.15001, 44.53999, 45.94, 47.32, 48.71001, 50.14001, 
    51.60999, 53.09001, 54.57, 56.07, 57.62, 59.21998, 60.83, 62.46998, 
    64.17001 ;

 Latitude =
  62.49, 62.91, 63.3, 63.65, 63.97, 64.26, 64.52, 64.77, 65.01, 65.23, 65.43, 
    65.62, 65.8, 65.98, 66.14, 66.3, 66.44, 66.58, 66.72, 66.85, 66.97, 
    67.09, 67.21, 67.32, 67.42, 67.53, 67.62, 67.72, 67.82, 67.91, 68, 68.08, 
    68.17, 68.25, 68.33, 68.41, 68.48, 68.56, 68.64, 68.71, 68.78, 68.85, 
    68.92, 68.98, 69.05, 69.11, 69.18, 69.24, 69.31, 69.37, 69.43, 69.49, 
    69.55, 69.61, 69.67, 69.73, 69.79, 69.84, 69.9, 69.96, 70.01, 70.07, 
    70.13, 70.18, 70.24, 70.29, 70.35, 70.4, 70.45, 70.51, 70.56, 70.61, 
    70.66, 70.72, 70.77, 70.82, 70.87, 70.92, 70.97, 71.01, 71.06, 71.1, 
    71.15, 71.19, 71.23, 71.26, 71.3, 71.33, 71.35, 71.37, 71.38, 71.38, 
    71.38, 71.35, 71.32, 71.26,
  62.59, 63.03, 63.41, 63.76, 64.08, 64.37, 64.64, 64.89, 65.13, 65.34, 
    65.55, 65.75, 65.93, 66.1, 66.26, 66.42, 66.57, 66.71, 66.85, 66.97, 
    67.1, 67.22, 67.34, 67.45, 67.55, 67.66, 67.76, 67.86, 67.95, 68.04, 
    68.13, 68.22, 68.3, 68.38, 68.46, 68.54, 68.62, 68.7, 68.77, 68.84, 
    68.92, 68.99, 69.06, 69.12, 69.19, 69.26, 69.32, 69.38, 69.45, 69.51, 
    69.57, 69.63, 69.7, 69.75, 69.81, 69.87, 69.93, 69.99, 70.05, 70.1, 
    70.16, 70.22, 70.27, 70.33, 70.38, 70.44, 70.5, 70.55, 70.6, 70.66, 
    70.71, 70.76, 70.82, 70.87, 70.92, 70.97, 71.02, 71.07, 71.12, 71.17, 
    71.21, 71.26, 71.3, 71.34, 71.38, 71.42, 71.45, 71.48, 71.51, 71.52, 
    71.54, 71.54, 71.53, 71.51, 71.47, 71.41,
  62.7, 63.14, 63.52, 63.87, 64.19, 64.49, 64.76, 65.01, 65.24, 65.47, 65.67, 
    65.87, 66.05, 66.22, 66.39, 66.55, 66.69, 66.83, 66.97, 67.1, 67.23, 
    67.35, 67.46, 67.57, 67.68, 67.79, 67.89, 67.99, 68.08, 68.18, 68.27, 
    68.35, 68.44, 68.52, 68.6, 68.68, 68.76, 68.83, 68.91, 68.98, 69.06, 
    69.13, 69.19, 69.26, 69.33, 69.4, 69.46, 69.53, 69.59, 69.65, 69.72, 
    69.78, 69.84, 69.9, 69.96, 70.02, 70.08, 70.14, 70.19, 70.25, 70.31, 
    70.36, 70.42, 70.48, 70.53, 70.59, 70.64, 70.7, 70.75, 70.81, 70.86, 
    70.91, 70.97, 71.02, 71.07, 71.12, 71.17, 71.22, 71.27, 71.32, 71.37, 
    71.41, 71.46, 71.5, 71.54, 71.57, 71.61, 71.64, 71.66, 71.68, 71.69, 
    71.69, 71.69, 71.66, 71.62, 71.56,
  62.8, 63.23, 63.63, 63.98, 64.3, 64.6, 64.87, 65.12, 65.36, 65.58, 65.79, 
    65.98, 66.17, 66.35, 66.51, 66.67, 66.82, 66.96, 67.1, 67.23, 67.35, 
    67.47, 67.59, 67.71, 67.81, 67.92, 68.02, 68.12, 68.22, 68.31, 68.4, 
    68.49, 68.57, 68.66, 68.74, 68.82, 68.9, 68.97, 69.05, 69.12, 69.19, 
    69.26, 69.33, 69.4, 69.47, 69.54, 69.6, 69.67, 69.73, 69.8, 69.86, 69.92, 
    69.98, 70.04, 70.1, 70.16, 70.22, 70.28, 70.34, 70.4, 70.45, 70.51, 
    70.57, 70.63, 70.68, 70.74, 70.79, 70.85, 70.9, 70.96, 71.01, 71.06, 
    71.12, 71.17, 71.22, 71.27, 71.33, 71.38, 71.43, 71.47, 71.52, 71.57, 
    71.61, 71.65, 71.69, 71.73, 71.76, 71.79, 71.82, 71.84, 71.85, 71.85, 
    71.84, 71.82, 71.78, 71.72,
  62.91, 63.35, 63.74, 64.09, 64.41, 64.71, 64.99, 65.24, 65.48, 65.7, 65.91, 
    66.11, 66.29, 66.47, 66.63, 66.79, 66.94, 67.09, 67.22, 67.35, 67.48, 
    67.6, 67.72, 67.83, 67.94, 68.05, 68.15, 68.25, 68.35, 68.44, 68.53, 
    68.62, 68.71, 68.79, 68.87, 68.95, 69.03, 69.11, 69.18, 69.26, 69.33, 
    69.4, 69.47, 69.54, 69.61, 69.68, 69.74, 69.81, 69.87, 69.94, 70, 70.06, 
    70.13, 70.19, 70.25, 70.31, 70.37, 70.43, 70.48, 70.54, 70.6, 70.66, 
    70.72, 70.77, 70.83, 70.89, 70.94, 71, 71.05, 71.11, 71.16, 71.22, 71.27, 
    71.32, 71.37, 71.43, 71.48, 71.53, 71.58, 71.63, 71.68, 71.72, 71.77, 
    71.81, 71.85, 71.88, 71.92, 71.95, 71.97, 71.99, 72, 72, 71.99, 71.97, 
    71.93, 71.87,
  63.02, 63.46, 63.85, 64.2, 64.53, 64.83, 65.1, 65.35, 65.59, 65.82, 66.03, 
    66.23, 66.41, 66.59, 66.76, 66.92, 67.07, 67.21, 67.35, 67.48, 67.61, 
    67.73, 67.85, 67.96, 68.07, 68.18, 68.28, 68.38, 68.48, 68.57, 68.67, 
    68.75, 68.84, 68.92, 69.01, 69.09, 69.17, 69.24, 69.32, 69.4, 69.47, 
    69.54, 69.61, 69.68, 69.75, 69.82, 69.88, 69.95, 70.01, 70.08, 70.14, 
    70.21, 70.27, 70.33, 70.39, 70.45, 70.51, 70.57, 70.63, 70.69, 70.75, 
    70.81, 70.86, 70.92, 70.98, 71.03, 71.09, 71.15, 71.2, 71.26, 71.31, 
    71.37, 71.42, 71.47, 71.53, 71.58, 71.63, 71.68, 71.73, 71.78, 71.83, 
    71.87, 71.92, 71.96, 72, 72.04, 72.07, 72.1, 72.13, 72.15, 72.16, 72.16, 
    72.15, 72.13, 72.08, 72.02,
  63.12, 63.56, 63.95, 64.31, 64.64, 64.93, 65.21, 65.47, 65.71, 65.93, 
    66.14, 66.34, 66.53, 66.71, 66.88, 67.04, 67.19, 67.33, 67.47, 67.61, 
    67.73, 67.86, 67.98, 68.09, 68.2, 68.31, 68.41, 68.51, 68.61, 68.7, 68.8, 
    68.89, 68.97, 69.06, 69.14, 69.22, 69.3, 69.38, 69.46, 69.53, 69.61, 
    69.68, 69.75, 69.82, 69.89, 69.96, 70.02, 70.09, 70.16, 70.22, 70.28, 
    70.35, 70.41, 70.47, 70.53, 70.6, 70.66, 70.72, 70.78, 70.83, 70.89, 
    70.95, 71.01, 71.07, 71.13, 71.18, 71.24, 71.3, 71.35, 71.41, 71.46, 
    71.52, 71.57, 71.63, 71.68, 71.73, 71.78, 71.84, 71.89, 71.93, 71.98, 
    72.03, 72.07, 72.12, 72.16, 72.19, 72.23, 72.26, 72.28, 72.3, 72.31, 
    72.31, 72.3, 72.28, 72.24, 72.17,
  63.22, 63.67, 64.07, 64.42, 64.75, 65.05, 65.33, 65.59, 65.82, 66.05, 
    66.26, 66.46, 66.65, 66.83, 67, 67.16, 67.31, 67.46, 67.6, 67.73, 67.86, 
    67.99, 68.11, 68.22, 68.33, 68.44, 68.54, 68.64, 68.74, 68.84, 68.93, 
    69.02, 69.11, 69.19, 69.28, 69.36, 69.44, 69.52, 69.59, 69.67, 69.74, 
    69.82, 69.89, 69.96, 70.03, 70.1, 70.16, 70.23, 70.3, 70.36, 70.43, 
    70.49, 70.55, 70.62, 70.68, 70.74, 70.8, 70.86, 70.92, 70.98, 71.04, 
    71.1, 71.16, 71.22, 71.27, 71.33, 71.39, 71.44, 71.5, 71.56, 71.61, 
    71.67, 71.72, 71.78, 71.83, 71.88, 71.94, 71.99, 72.04, 72.09, 72.14, 
    72.18, 72.23, 72.27, 72.31, 72.35, 72.38, 72.41, 72.44, 72.46, 72.47, 
    72.47, 72.46, 72.44, 72.39, 72.33,
  63.33, 63.77, 64.17, 64.53, 64.86, 65.16, 65.44, 65.7, 65.94, 66.17, 66.38, 
    66.58, 66.77, 66.95, 67.12, 67.28, 67.43, 67.58, 67.72, 67.86, 67.99, 
    68.11, 68.23, 68.35, 68.46, 68.57, 68.67, 68.77, 68.87, 68.97, 69.06, 
    69.15, 69.24, 69.33, 69.41, 69.49, 69.57, 69.65, 69.73, 69.81, 69.88, 
    69.95, 70.03, 70.1, 70.17, 70.24, 70.3, 70.37, 70.44, 70.5, 70.57, 70.63, 
    70.7, 70.76, 70.82, 70.88, 70.94, 71.01, 71.07, 71.13, 71.19, 71.24, 
    71.3, 71.36, 71.42, 71.48, 71.54, 71.59, 71.65, 71.71, 71.76, 71.82, 
    71.87, 71.93, 71.98, 72.03, 72.09, 72.14, 72.19, 72.24, 72.29, 72.34, 
    72.38, 72.43, 72.47, 72.5, 72.54, 72.57, 72.59, 72.61, 72.62, 72.62, 
    72.61, 72.59, 72.55, 72.48,
  63.42, 63.87, 64.28, 64.64, 64.97, 65.27, 65.55, 65.81, 66.05, 66.28, 
    66.49, 66.7, 66.89, 67.07, 67.24, 67.4, 67.56, 67.71, 67.85, 67.98, 
    68.11, 68.24, 68.36, 68.47, 68.59, 68.69, 68.8, 68.9, 69, 69.1, 69.19, 
    69.28, 69.37, 69.46, 69.54, 69.63, 69.71, 69.79, 69.87, 69.94, 70.02, 
    70.09, 70.16, 70.24, 70.31, 70.37, 70.44, 70.51, 70.58, 70.64, 70.71, 
    70.78, 70.84, 70.9, 70.96, 71.03, 71.09, 71.15, 71.21, 71.27, 71.33, 
    71.39, 71.45, 71.51, 71.57, 71.63, 71.68, 71.74, 71.8, 71.86, 71.91, 
    71.97, 72.02, 72.08, 72.13, 72.19, 72.24, 72.29, 72.34, 72.39, 72.44, 
    72.49, 72.54, 72.58, 72.62, 72.66, 72.69, 72.72, 72.75, 72.77, 72.78, 
    72.78, 72.77, 72.74, 72.7, 72.63,
  63.54, 63.99, 64.38, 64.74, 65.08, 65.38, 65.67, 65.92, 66.17, 66.4, 66.61, 
    66.82, 67.01, 67.19, 67.36, 67.52, 67.68, 67.83, 67.97, 68.1, 68.24, 
    68.36, 68.48, 68.6, 68.71, 68.82, 68.93, 69.03, 69.13, 69.23, 69.32, 
    69.42, 69.5, 69.59, 69.68, 69.76, 69.84, 69.92, 70, 70.08, 70.15, 70.23, 
    70.3, 70.37, 70.44, 70.51, 70.58, 70.65, 70.72, 70.79, 70.85, 70.92, 
    70.98, 71.04, 71.11, 71.17, 71.23, 71.29, 71.36, 71.42, 71.48, 71.54, 
    71.6, 71.66, 71.72, 71.77, 71.83, 71.89, 71.95, 72.01, 72.06, 72.12, 
    72.17, 72.23, 72.28, 72.34, 72.39, 72.45, 72.5, 72.55, 72.6, 72.65, 
    72.69, 72.74, 72.78, 72.82, 72.85, 72.88, 72.9, 72.92, 72.93, 72.93, 
    72.92, 72.9, 72.85, 72.78,
  63.63, 64.08, 64.48, 64.85, 65.19, 65.49, 65.77, 66.03, 66.28, 66.51, 
    66.73, 66.93, 67.12, 67.31, 67.48, 67.64, 67.8, 67.95, 68.09, 68.23, 
    68.36, 68.49, 68.61, 68.73, 68.84, 68.95, 69.06, 69.16, 69.26, 69.36, 
    69.45, 69.55, 69.64, 69.72, 69.81, 69.89, 69.98, 70.06, 70.14, 70.21, 
    70.29, 70.36, 70.44, 70.51, 70.58, 70.65, 70.72, 70.79, 70.86, 70.93, 
    70.99, 71.06, 71.12, 71.19, 71.25, 71.31, 71.38, 71.44, 71.5, 71.56, 
    71.62, 71.68, 71.74, 71.8, 71.86, 71.92, 71.98, 72.04, 72.1, 72.15, 
    72.21, 72.27, 72.32, 72.38, 72.44, 72.49, 72.54, 72.6, 72.65, 72.7, 
    72.75, 72.8, 72.85, 72.89, 72.93, 72.97, 73, 73.04, 73.06, 73.08, 73.09, 
    73.09, 73.08, 73.05, 73.01, 72.94 ;

 Longitude =
  132.83, 133.74, 134.6, 135.4, 136.16, 136.87, 137.55, 138.21, 138.85, 
    139.46, 140.03, 140.59, 141.14, 141.67, 142.19, 142.69, 143.17, 143.64, 
    144.11, 144.57, 145, 145.44, 145.87, 146.29, 146.71, 147.11, 147.5, 
    147.9, 148.3, 148.69, 149.06, 149.44, 149.82, 150.19, 150.56, 150.93, 
    151.3, 151.66, 152.03, 152.39, 152.75, 153.11, 153.48, 153.85, 154.21, 
    154.57, 154.93, 155.3, 155.68, 156.05, 156.42, 156.8, 157.18, 157.57, 
    157.96, 158.35, 158.75, 159.16, 159.57, 159.98, 160.4, 160.83, 161.27, 
    161.73, 162.18, 162.64, 163.11, 163.61, 164.11, 164.62, 165.14, 165.68, 
    166.24, 166.82, 167.41, 168.01, 168.66, 169.32, 170.02, 170.72, 171.45, 
    172.22, 173.05, 173.91, 174.79, 175.72, 176.72, 177.77, 178.89, -179.93, 
    -178.67, -177.31, -175.84, -174.25, -172.55, -170.69,
  132.58, 133.5, 134.35, 135.15, 135.9, 136.62, 137.31, 137.97, 138.59, 
    139.19, 139.78, 140.35, 140.9, 141.43, 141.93, 142.43, 142.93, 143.41, 
    143.87, 144.31, 144.76, 145.2, 145.63, 146.05, 146.46, 146.87, 147.27, 
    147.67, 148.06, 148.45, 148.83, 149.22, 149.59, 149.96, 150.33, 150.71, 
    151.08, 151.45, 151.81, 152.17, 152.54, 152.9, 153.27, 153.63, 153.99, 
    154.36, 154.73, 155.1, 155.47, 155.85, 156.23, 156.61, 156.99, 157.38, 
    157.77, 158.16, 158.57, 158.98, 159.38, 159.8, 160.23, 160.66, 161.11, 
    161.55, 162.01, 162.48, 162.96, 163.45, 163.95, 164.47, 165, 165.55, 
    166.11, 166.68, 167.27, 167.9, 168.55, 169.21, 169.89, 170.61, 171.36, 
    172.15, 172.96, 173.81, 174.72, 175.67, 176.67, 177.73, 178.83, -179.97, 
    -178.67, -177.29, -175.83, -174.25, -172.53, -170.62,
  132.34, 133.25, 134.09, 134.89, 135.65, 136.37, 137.06, 137.71, 138.34, 
    138.95, 139.54, 140.1, 140.64, 141.17, 141.69, 142.19, 142.68, 143.15, 
    143.61, 144.07, 144.52, 144.96, 145.38, 145.81, 146.22, 146.64, 147.04, 
    147.43, 147.82, 148.22, 148.61, 148.98, 149.36, 149.73, 150.11, 150.49, 
    150.85, 151.22, 151.59, 151.96, 152.32, 152.69, 153.05, 153.42, 153.79, 
    154.16, 154.52, 154.89, 155.27, 155.65, 156.03, 156.41, 156.79, 157.18, 
    157.58, 157.98, 158.38, 158.79, 159.2, 159.63, 160.06, 160.48, 160.93, 
    161.38, 161.85, 162.32, 162.8, 163.29, 163.8, 164.33, 164.86, 165.4, 
    165.96, 166.55, 167.15, 167.78, 168.42, 169.09, 169.79, 170.52, 171.27, 
    172.05, 172.87, 173.74, 174.66, 175.6, 176.6, 177.66, 178.81, -179.97, 
    -178.68, -177.32, -175.84, -174.23, -172.47, -170.57,
  132.07, 132.97, 133.83, 134.64, 135.39, 136.1, 136.78, 137.45, 138.09, 
    138.69, 139.27, 139.83, 140.39, 140.92, 141.44, 141.94, 142.42, 142.9, 
    143.37, 143.83, 144.27, 144.7, 145.14, 145.57, 145.98, 146.39, 146.79, 
    147.2, 147.59, 147.98, 148.37, 148.75, 149.13, 149.51, 149.88, 150.25, 
    150.63, 151, 151.37, 151.73, 152.1, 152.46, 152.84, 153.21, 153.57, 
    153.94, 154.31, 154.69, 155.07, 155.44, 155.82, 156.21, 156.6, 156.99, 
    157.39, 157.78, 158.19, 158.61, 159.02, 159.44, 159.87, 160.31, 160.76, 
    161.22, 161.68, 162.15, 162.64, 163.14, 163.65, 164.17, 164.7, 165.26, 
    165.83, 166.42, 167.02, 167.64, 168.3, 168.99, 169.69, 170.4, 171.16, 
    171.95, 172.79, 173.67, 174.57, 175.53, 176.55, 177.64, 178.78, 179.98, 
    -178.72, -177.31, -175.8, -174.19, -172.46, -170.55,
  131.82, 132.73, 133.58, 134.37, 135.13, 135.85, 136.54, 137.2, 137.82, 
    138.43, 139.02, 139.59, 140.14, 140.66, 141.17, 141.68, 142.18, 142.66, 
    143.12, 143.57, 144.02, 144.46, 144.9, 145.32, 145.73, 146.15, 146.56, 
    146.96, 147.35, 147.74, 148.13, 148.52, 148.9, 149.27, 149.64, 150.02, 
    150.4, 150.77, 151.14, 151.5, 151.88, 152.25, 152.62, 152.98, 153.35, 
    153.73, 154.11, 154.48, 154.85, 155.23, 155.62, 156.01, 156.4, 156.79, 
    157.19, 157.59, 158, 158.42, 158.83, 159.26, 159.69, 160.14, 160.58, 
    161.04, 161.51, 161.99, 162.48, 162.98, 163.49, 164.02, 164.56, 165.12, 
    165.69, 166.27, 166.88, 167.53, 168.19, 168.86, 169.56, 170.29, 171.07, 
    171.87, 172.7, 173.57, 174.5, 175.49, 176.51, 177.58, 178.72, 179.96, 
    -178.71, -177.3, -175.82, -174.2, -172.42, -170.46,
  131.57, 132.47, 133.31, 134.11, 134.87, 135.59, 136.27, 136.92, 137.56, 
    138.17, 138.76, 139.32, 139.86, 140.4, 140.92, 141.43, 141.92, 142.39, 
    142.86, 143.32, 143.77, 144.21, 144.64, 145.07, 145.49, 145.9, 146.31, 
    146.71, 147.11, 147.5, 147.89, 148.27, 148.65, 149.03, 149.42, 149.79, 
    150.16, 150.54, 150.91, 151.28, 151.65, 152.02, 152.39, 152.77, 153.14, 
    153.51, 153.88, 154.26, 154.65, 155.03, 155.42, 155.8, 156.19, 156.59, 
    157, 157.4, 157.8, 158.22, 158.64, 159.08, 159.51, 159.95, 160.4, 160.87, 
    161.34, 161.82, 162.31, 162.81, 163.33, 163.87, 164.41, 164.96, 165.54, 
    166.14, 166.76, 167.39, 168.05, 168.74, 169.45, 170.2, 170.96, 171.76, 
    172.61, 173.5, 174.44, 175.4, 176.43, 177.53, 178.7, 179.95, -178.75, 
    -177.34, -175.81, -174.16, -172.36, -170.43,
  131.29, 132.19, 133.05, 133.85, 134.6, 135.31, 136, 136.66, 137.3, 137.9, 
    138.49, 139.05, 139.61, 140.15, 140.66, 141.16, 141.65, 142.14, 142.61, 
    143.06, 143.51, 143.95, 144.39, 144.82, 145.24, 145.65, 146.06, 146.46, 
    146.86, 147.25, 147.64, 148.03, 148.42, 148.8, 149.17, 149.55, 149.93, 
    150.31, 150.68, 151.05, 151.42, 151.79, 152.17, 152.55, 152.92, 153.29, 
    153.67, 154.05, 154.43, 154.81, 155.2, 155.59, 155.99, 156.39, 156.79, 
    157.19, 157.61, 158.03, 158.46, 158.88, 159.32, 159.77, 160.23, 160.69, 
    161.16, 161.64, 162.14, 162.65, 163.17, 163.7, 164.25, 164.82, 165.41, 
    166, 166.61, 167.25, 167.93, 168.63, 169.34, 170.08, 170.85, 171.67, 
    172.53, 173.42, 174.35, 175.33, 176.38, 177.49, 178.66, 179.89, -178.78, 
    -177.33, -175.79, -174.14, -172.36, -170.39,
  131.03, 131.94, 132.79, 133.58, 134.33, 135.05, 135.74, 136.4, 137.03, 
    137.63, 138.23, 138.8, 139.35, 139.87, 140.39, 140.9, 141.4, 141.88, 
    142.34, 142.8, 143.25, 143.7, 144.14, 144.56, 144.98, 145.4, 145.81, 
    146.21, 146.61, 147, 147.4, 147.79, 148.17, 148.55, 148.93, 149.32, 
    149.7, 150.07, 150.44, 150.81, 151.19, 151.57, 151.94, 152.31, 152.69, 
    153.07, 153.45, 153.83, 154.21, 154.6, 154.99, 155.39, 155.78, 156.17, 
    156.58, 157, 157.42, 157.83, 158.25, 158.69, 159.13, 159.59, 160.04, 
    160.51, 160.99, 161.48, 161.98, 162.48, 163, 163.54, 164.1, 164.67, 
    165.25, 165.85, 166.48, 167.13, 167.8, 168.49, 169.21, 169.97, 170.76, 
    171.58, 172.42, 173.32, 174.28, 175.28, 176.32, 177.42, 178.6, 179.88, 
    -178.76, -177.32, -175.8, -174.14, -172.31, -170.3,
  130.77, 131.67, 132.51, 133.31, 134.07, 134.79, 135.47, 136.12, 136.76, 
    137.38, 137.96, 138.52, 139.07, 139.61, 140.14, 140.64, 141.13, 141.61, 
    142.08, 142.54, 142.99, 143.43, 143.87, 144.3, 144.73, 145.14, 145.55, 
    145.95, 146.36, 146.76, 147.15, 147.53, 147.92, 148.31, 148.69, 149.07, 
    149.45, 149.83, 150.21, 150.58, 150.96, 151.33, 151.71, 152.09, 152.47, 
    152.84, 153.22, 153.6, 154, 154.39, 154.78, 155.17, 155.56, 155.97, 
    156.38, 156.79, 157.2, 157.63, 158.06, 158.5, 158.94, 159.39, 159.85, 
    160.33, 160.81, 161.3, 161.79, 162.31, 162.84, 163.39, 163.94, 164.51, 
    165.1, 165.71, 166.34, 166.99, 167.66, 168.37, 169.11, 169.87, 170.65, 
    171.46, 172.34, 173.25, 174.21, 175.2, 176.25, 177.38, 178.58, 179.85, 
    -178.8, -177.36, -175.79, -174.09, -172.26, -170.28,
  130.49, 131.39, 132.25, 133.04, 133.79, 134.5, 135.19, 135.86, 136.49, 
    137.09, 137.68, 138.25, 138.81, 139.35, 139.86, 140.36, 140.86, 141.35, 
    141.82, 142.27, 142.72, 143.17, 143.62, 144.05, 144.46, 144.88, 145.29, 
    145.71, 146.11, 146.5, 146.89, 147.29, 147.68, 148.06, 148.44, 148.82, 
    149.21, 149.59, 149.97, 150.34, 150.71, 151.1, 151.48, 151.86, 152.23, 
    152.61, 153, 153.39, 153.77, 154.16, 154.55, 154.96, 155.36, 155.76, 
    156.16, 156.58, 157.01, 157.43, 157.86, 158.29, 158.74, 159.2, 159.67, 
    160.14, 160.62, 161.12, 161.63, 162.15, 162.67, 163.21, 163.78, 164.36, 
    164.96, 165.56, 166.19, 166.85, 167.54, 168.25, 168.98, 169.73, 170.53, 
    171.38, 172.25, 173.16, 174.11, 175.13, 176.21, 177.34, 178.53, 179.81, 
    -178.82, -177.33, -175.76, -174.08, -172.25, -170.22,
  130.23, 131.14, 131.97, 132.76, 133.52, 134.24, 134.93, 135.58, 136.21, 
    136.82, 137.42, 137.99, 138.53, 139.06, 139.59, 140.1, 140.6, 141.08, 
    141.54, 142.01, 142.46, 142.91, 143.35, 143.78, 144.2, 144.62, 145.04, 
    145.44, 145.84, 146.25, 146.65, 147.04, 147.42, 147.8, 148.19, 148.58, 
    148.97, 149.34, 149.72, 150.1, 150.48, 150.86, 151.24, 151.62, 152, 
    152.39, 152.77, 153.15, 153.54, 153.94, 154.34, 154.74, 155.13, 155.54, 
    155.96, 156.38, 156.8, 157.22, 157.65, 158.1, 158.55, 159.01, 159.47, 
    159.95, 160.44, 160.94, 161.45, 161.96, 162.5, 163.06, 163.62, 164.2, 
    164.79, 165.41, 166.05, 166.72, 167.4, 168.11, 168.85, 169.63, 170.44, 
    171.27, 172.14, 173.07, 174.05, 175.07, 176.14, 177.26, 178.49, 179.8, 
    -178.82, -177.35, -175.77, -174.05, -172.17, -170.13,
  129.95, 130.85, 131.69, 132.49, 133.25, 133.96, 134.64, 135.3, 135.94, 
    136.55, 137.14, 137.7, 138.25, 138.8, 139.32, 139.82, 140.32, 140.8, 
    141.28, 141.74, 142.19, 142.64, 143.08, 143.52, 143.94, 144.36, 144.77, 
    145.18, 145.59, 145.99, 146.38, 146.77, 147.17, 147.56, 147.94, 148.33, 
    148.71, 149.09, 149.48, 149.86, 150.23, 150.61, 151, 151.39, 151.77, 
    152.15, 152.53, 152.92, 153.32, 153.72, 154.11, 154.51, 154.92, 155.33, 
    155.74, 156.16, 156.58, 157.02, 157.46, 157.9, 158.35, 158.81, 159.28, 
    159.77, 160.26, 160.75, 161.26, 161.79, 162.34, 162.89, 163.45, 164.03, 
    164.64, 165.27, 165.91, 166.57, 167.26, 167.99, 168.74, 169.51, 170.31, 
    171.16, 172.06, 173, 173.96, 174.98, 176.07, 177.24, 178.46, 179.76, 
    -178.86, -177.36, -175.74, -174.01, -172.14, -170.12 ;

 Orb_mode = 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 Polo = 2, 2, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 2, 3, 3, 3, 3, 3, 3 ;

 PrecipType =
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888 ;

 Prob_SF =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 33, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 65, 66, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 42, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 66, 65, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 61, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 57, 49, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 56, 55, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 57, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 49, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 44, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 53, 53, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 64, 64, 
    56, 63, 62, 61, 64, 61, 59, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 64, 0, 62, 64, 
    65, 64, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 Qc =
  1, 0, 144, 8192,
  1, 0, 144, 8192,
  1, 0, 144, 8192,
  1, 0, 144, 8192,
  1, 0, 144, 8192,
  0, 0, 128, 8192,
  0, 0, 128, 8192,
  0, 0, 128, 8192,
  1, 0, 132, 8192,
  1, 0, 188, 8192,
  1, 12, 3776, 8192,
  1, 12, 3788, 8192,
  1, 12, 3788, 8192,
  1, 12, 3804, 8192,
  1, 0, 172, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 172, 8192,
  0, 0, 160, 8192,
  0, 0, 160, 8192,
  0, 0, 160, 8192,
  1, 0, 164, 8192,
  1, 0, 176, 8192,
  1, 0, 188, 8192,
  1, 0, 164, 8192,
  1, 0, 164, 8192,
  1, 0, 188, 8192,
  1, 0, 180, 8192,
  1, 0, 180, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 180, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 180, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 176, 8192,
  1, 0, 176, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 156, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 12, 3776, 8192,
  1, 0, 156, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 176, 8192,
  1, 0, 176, 8192,
  1, 0, 176, 8192,
  1, 0, 180, 8192,
  1, 0, 188, 8192,
  1, 0, 180, 8192,
  0, 0, 128, 0,
  1, 0, 144, 0,
  1, 0, 16, 4096,
  1, 0, 48, 4096,
  1, 0, 48, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 48, 4096,
  1, 0, 48, 4096,
  1, 0, 20, 4096,
  1, 0, 48, 4096,
  1, 0, 48, 4096,
  1, 0, 48, 4096,
  0, 0, 32, 4096,
  1, 0, 144, 0,
  1, 0, 144, 0,
  0, 0, 0, 4096,
  0, 0, 160, 8192,
  0, 0, 160, 8192,
  1, 0, 144, 0,
  1, 0, 144, 0,
  1, 0, 144, 0,
  1, 0, 144, 0,
  1, 0, 144, 0,
  1, 0, 144, 8192,
  1, 0, 144, 8192,
  1, 0, 144, 8192,
  1, 0, 148, 8192,
  0, 0, 128, 8192,
  0, 0, 128, 8192,
  0, 0, 128, 8192,
  1, 0, 172, 8192,
  1, 0, 172, 8192,
  1, 12, 3776, 8192,
  1, 12, 3788, 8192,
  1, 12, 3788, 8192,
  1, 12, 3776, 8192,
  1, 12, 3776, 8192,
  1, 0, 172, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 172, 8192,
  0, 0, 160, 8192,
  0, 0, 160, 8192,
  0, 0, 160, 8192,
  1, 0, 180, 8192,
  1, 0, 180, 8192,
  1, 0, 188, 8192,
  1, 0, 176, 8192,
  1, 0, 180, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 164, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 156, 8192,
  1, 0, 172, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 176, 8192,
  1, 0, 176, 8192,
  1, 0, 188, 8192,
  1, 0, 176, 8192,
  1, 0, 176, 8192,
  1, 0, 176, 8192,
  1, 0, 180, 8192,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 48, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 52, 4096,
  1, 0, 48, 4096,
  1, 0, 20, 4096,
  1, 0, 52, 4096,
  1, 0, 48, 4096,
  1, 0, 48, 4096,
  0, 0, 32, 4096,
  0, 0, 0, 4096,
  1, 0, 144, 0,
  0, 0, 32, 4096,
  0, 0, 32, 4096,
  1, 0, 144, 0,
  1, 0, 144, 0,
  1, 0, 144, 0,
  1, 0, 144, 0,
  1, 0, 144, 0,
  1, 0, 144, 0,
  1, 0, 144, 8192,
  1, 0, 144, 8192,
  1, 0, 144, 8192,
  0, 0, 128, 8192,
  0, 0, 128, 8192,
  0, 0, 128, 8192,
  1, 0, 132, 8192,
  1, 0, 172, 8192,
  1, 12, 3776, 8192,
  1, 12, 3788, 8192,
  1, 12, 3776, 8192,
  1, 12, 3776, 8192,
  1, 12, 3776, 8192,
  1, 0, 172, 8192,
  1, 0, 188, 8192,
  1, 0, 172, 8192,
  1, 0, 188, 8192,
  1, 0, 172, 8192,
  0, 0, 160, 8192,
  0, 0, 160, 8192,
  1, 0, 180, 8192,
  1, 0, 164, 8192,
  1, 0, 176, 8192,
  1, 0, 176, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 172, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 176, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 180, 8192,
  1, 0, 180, 8192,
  1, 0, 188, 8192,
  0, 0, 160, 8192,
  1, 0, 188, 8192,
  1, 0, 156, 8192,
  1, 0, 172, 8192,
  1, 0, 176, 8192,
  1, 0, 176, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 176, 8192,
  1, 0, 144, 8192,
  1, 0, 176, 8192,
  1, 0, 176, 8192,
  1, 0, 176, 8192,
  1, 0, 176, 8192,
  1, 0, 16, 4096,
  1, 0, 20, 4096,
  1, 0, 48, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 48, 4096,
  1, 0, 48, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 20, 4096,
  1, 0, 20, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 48, 4096,
  0, 0, 32, 4096,
  0, 0, 0, 4096,
  0, 0, 0, 4096,
  0, 0, 0, 4096,
  1, 0, 144, 0,
  0, 0, 0, 4096,
  1, 0, 144, 0,
  1, 0, 144, 0,
  1, 0, 144, 0,
  1, 0, 144, 0,
  1, 0, 144, 0,
  1, 0, 144, 0,
  1, 0, 144, 8192,
  0, 0, 128, 8192,
  0, 0, 128, 8192,
  0, 0, 128, 8192,
  0, 0, 128, 8192,
  0, 0, 128, 8192,
  1, 0, 172, 8192,
  0, 0, 160, 8192,
  1, 12, 3776, 8192,
  1, 12, 3788, 8192,
  1, 12, 3776, 8192,
  1, 12, 3776, 8192,
  0, 0, 160, 8192,
  1, 0, 188, 8192,
  1, 0, 172, 8192,
  1, 0, 172, 8192,
  1, 0, 188, 8192,
  1, 0, 172, 8192,
  1, 0, 172, 8192,
  0, 0, 160, 8192,
  0, 0, 160, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 164, 8192,
  1, 0, 176, 8192,
  0, 0, 160, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 176, 8192,
  1, 0, 180, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  0, 0, 160, 8192,
  1, 0, 176, 8192,
  1, 0, 176, 8192,
  1, 0, 180, 8192,
  1, 0, 188, 8192,
  1, 0, 176, 8192,
  1, 0, 176, 8192,
  1, 0, 176, 8192,
  1, 0, 176, 8192,
  1, 0, 176, 8192,
  1, 0, 176, 8192,
  1, 0, 176, 8192,
  0, 0, 0, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 48, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 48, 4096,
  1, 0, 48, 4096,
  1, 0, 48, 4096,
  1, 0, 16, 4096,
  1, 0, 20, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  0, 0, 0, 4096,
  1, 0, 48, 4096,
  1, 0, 48, 4096,
  0, 0, 32, 4096,
  0, 0, 0, 4096,
  0, 0, 0, 4096,
  0, 0, 0, 4096,
  0, 0, 32, 4096,
  1, 0, 144, 0,
  1, 0, 144, 0,
  0, 0, 128, 0,
  1, 0, 144, 0,
  1, 0, 144, 0,
  1, 0, 144, 0,
  0, 0, 128, 8192,
  0, 0, 128, 8192,
  0, 0, 128, 8192,
  0, 0, 128, 8192,
  0, 0, 128, 8192,
  0, 0, 160, 8192,
  1, 0, 172, 8192,
  0, 0, 160, 8192,
  1, 12, 3776, 8192,
  1, 12, 3776, 8192,
  1, 12, 3776, 8192,
  1, 12, 3776, 8192,
  0, 0, 160, 8192,
  1, 0, 172, 8192,
  0, 0, 160, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 172, 8192,
  1, 0, 188, 8192,
  1, 0, 164, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 176, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 172, 8192,
  1, 0, 180, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 180, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 180, 8192,
  1, 0, 176, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 176, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 176, 8192,
  1, 0, 176, 8192,
  1, 0, 176, 8192,
  1, 0, 176, 8192,
  1, 0, 176, 8192,
  1, 0, 176, 8192,
  1, 0, 176, 8192,
  1, 0, 176, 8192,
  0, 0, 0, 4096,
  1, 0, 144, 8192,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 48, 4096,
  1, 0, 48, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 20, 4096,
  1, 0, 16, 4096,
  1, 0, 48, 4096,
  1, 0, 48, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 20, 4096,
  0, 0, 128, 0,
  0, 0, 128, 0,
  1, 0, 144, 0,
  1, 0, 48, 4096,
  0, 0, 32, 4096,
  0, 0, 0, 4096,
  0, 0, 0, 4096,
  1, 0, 4, 4096,
  1, 0, 144, 0,
  1, 0, 144, 0,
  1, 0, 144, 0,
  1, 0, 144, 0,
  1, 0, 144, 0,
  0, 0, 128, 0,
  1, 0, 144, 0,
  0, 0, 128, 8192,
  0, 0, 160, 8192,
  0, 0, 160, 8192,
  0, 0, 128, 8192,
  0, 0, 160, 8192,
  0, 0, 128, 8192,
  0, 0, 160, 8192,
  1, 12, 3776, 8192,
  1, 12, 3776, 8192,
  1, 12, 3776, 8192,
  0, 0, 160, 8192,
  1, 0, 172, 8192,
  0, 0, 160, 8192,
  1, 0, 172, 8192,
  1, 0, 172, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 180, 8192,
  1, 0, 180, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 164, 8192,
  1, 0, 176, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 180, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 172, 8192,
  1, 0, 188, 8192,
  1, 0, 180, 8192,
  1, 0, 188, 8192,
  1, 0, 180, 8192,
  1, 0, 188, 8192,
  1, 0, 172, 8192,
  1, 0, 176, 8192,
  1, 0, 176, 8192,
  1, 0, 176, 8192,
  1, 0, 176, 8192,
  1, 0, 176, 8192,
  1, 0, 176, 8192,
  1, 0, 176, 8192,
  1, 0, 176, 8192,
  0, 0, 0, 4096,
  0, 0, 0, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 48, 4096,
  1, 0, 16, 4096,
  1, 0, 20, 4096,
  1, 0, 16, 4096,
  1, 0, 48, 4096,
  1, 0, 48, 4096,
  1, 0, 48, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 144, 0,
  1, 0, 144, 0,
  1, 0, 144, 0,
  1, 0, 48, 4096,
  0, 0, 32, 4096,
  0, 0, 0, 4096,
  0, 0, 0, 4096,
  0, 0, 0, 4096,
  1, 0, 144, 0,
  1, 0, 144, 0,
  1, 0, 144, 0,
  1, 0, 144, 0,
  1, 0, 144, 0,
  1, 0, 144, 0,
  1, 0, 148, 0,
  0, 0, 160, 8192,
  0, 0, 160, 8192,
  0, 0, 160, 8192,
  1, 0, 172, 8192,
  0, 0, 160, 8192,
  1, 0, 164, 8192,
  0, 0, 160, 8192,
  1, 12, 3776, 8192,
  1, 12, 3780, 8192,
  0, 0, 160, 8192,
  0, 0, 160, 8192,
  0, 0, 160, 8192,
  0, 0, 160, 8192,
  0, 0, 160, 8192,
  1, 0, 172, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 180, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 172, 8192,
  0, 0, 160, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 176, 8192,
  1, 0, 188, 8192,
  1, 0, 172, 8192,
  1, 0, 176, 8192,
  1, 0, 188, 8192,
  1, 0, 180, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 172, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 176, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  0, 0, 160, 8192,
  1, 0, 176, 8192,
  1, 0, 176, 8192,
  1, 0, 144, 8192,
  1, 0, 176, 8192,
  1, 0, 176, 8192,
  1, 0, 176, 8192,
  1, 0, 176, 8192,
  1, 0, 176, 8192,
  1, 0, 176, 8192,
  0, 0, 0, 4096,
  1, 0, 144, 0,
  0, 0, 0, 4096,
  1, 0, 16, 4096,
  1, 0, 48, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 48, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 20, 4096,
  1, 0, 16, 4096,
  1, 0, 48, 4096,
  1, 0, 48, 4096,
  1, 0, 48, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 48, 4096,
  1, 0, 144, 0,
  1, 0, 144, 0,
  1, 0, 48, 4096,
  1, 0, 48, 4096,
  0, 0, 0, 4096,
  0, 0, 0, 4096,
  0, 0, 0, 4096,
  0, 0, 0, 4096,
  1, 0, 144, 0,
  1, 0, 144, 0,
  1, 0, 144, 0,
  1, 0, 144, 0,
  1, 0, 148, 0,
  1, 0, 144, 0,
  1, 0, 144, 0,
  0, 0, 160, 8192,
  0, 0, 160, 8192,
  0, 0, 160, 8192,
  0, 0, 160, 8192,
  0, 0, 160, 8192,
  0, 0, 160, 8192,
  1, 12, 3776, 8192,
  1, 12, 3776, 8192,
  1, 12, 3776, 8192,
  1, 0, 172, 8192,
  1, 0, 172, 8192,
  1, 0, 172, 8192,
  0, 0, 160, 8192,
  0, 0, 160, 8192,
  0, 0, 160, 8192,
  1, 0, 180, 8192,
  1, 0, 180, 8192,
  0, 0, 160, 8192,
  1, 0, 180, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 176, 8192,
  1, 0, 180, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 176, 8192,
  1, 0, 176, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 172, 8192,
  1, 0, 172, 8192,
  0, 0, 160, 8192,
  1, 0, 172, 8192,
  1, 0, 188, 8192,
  1, 0, 172, 8192,
  1, 0, 172, 8192,
  1, 0, 172, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 172, 8192,
  1, 0, 172, 8192,
  1, 0, 188, 8192,
  1, 0, 176, 8192,
  1, 0, 188, 8192,
  1, 0, 172, 8192,
  1, 0, 176, 8192,
  0, 0, 160, 8192,
  0, 0, 160, 8192,
  1, 0, 176, 8192,
  1, 0, 176, 8192,
  1, 0, 176, 8192,
  1, 0, 176, 8192,
  1, 0, 176, 8192,
  1, 0, 176, 8192,
  1, 0, 176, 8192,
  1, 0, 144, 8192,
  1, 0, 16, 4096,
  0, 0, 0, 4096,
  1, 0, 16, 4096,
  1, 0, 48, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 20, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 20, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 28, 4096,
  1, 0, 28, 4096,
  1, 0, 48, 4096,
  1, 0, 48, 4096,
  1, 0, 48, 4096,
  1, 0, 48, 4096,
  1, 0, 16, 4096,
  1, 0, 48, 4096,
  1, 0, 48, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  0, 0, 0, 4096,
  0, 0, 0, 4096,
  0, 0, 0, 4096,
  0, 0, 0, 4096,
  0, 0, 0, 4096,
  1, 0, 144, 0,
  1, 0, 144, 0,
  1, 0, 144, 0,
  1, 0, 148, 0,
  1, 0, 156, 0,
  1, 0, 156, 0,
  1, 0, 144, 0,
  0, 0, 160, 8192,
  0, 0, 160, 8192,
  0, 0, 160, 8192,
  0, 0, 160, 8192,
  0, 0, 160, 8192,
  1, 12, 3776, 8192,
  1, 12, 3776, 8192,
  0, 0, 160, 8192,
  0, 0, 160, 8192,
  0, 0, 160, 8192,
  0, 0, 160, 8192,
  1, 0, 172, 8192,
  0, 0, 160, 8192,
  0, 0, 160, 8192,
  0, 0, 160, 8192,
  1, 0, 164, 8192,
  1, 0, 180, 8192,
  0, 0, 160, 8192,
  1, 0, 180, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 176, 8192,
  1, 0, 164, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 172, 8192,
  1, 0, 164, 8192,
  1, 0, 172, 8192,
  1, 0, 172, 8192,
  1, 0, 172, 8192,
  1, 0, 172, 8192,
  1, 0, 172, 8192,
  1, 0, 172, 8192,
  1, 0, 172, 8192,
  1, 0, 172, 8192,
  1, 0, 188, 8192,
  1, 0, 176, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 176, 8192,
  1, 0, 176, 8192,
  1, 0, 176, 8192,
  1, 0, 176, 8192,
  0, 0, 160, 8192,
  0, 0, 160, 8192,
  0, 0, 160, 8192,
  1, 0, 176, 8192,
  1, 0, 176, 8192,
  1, 0, 176, 8192,
  1, 0, 48, 4096,
  0, 0, 0, 4096,
  0, 0, 0, 4096,
  1, 0, 16, 4096,
  1, 0, 48, 4096,
  1, 0, 52, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 20, 4096,
  1, 0, 16, 4096,
  1, 0, 20, 4096,
  1, 0, 16, 4096,
  1, 0, 48, 4096,
  1, 0, 48, 4096,
  1, 0, 52, 4096,
  1, 0, 48, 4096,
  1, 0, 48, 4096,
  1, 0, 48, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  0, 0, 0, 4096,
  0, 0, 32, 4096,
  0, 0, 32, 4096,
  1, 0, 144, 0,
  1, 0, 144, 0,
  1, 0, 144, 0,
  1, 0, 144, 0,
  1, 0, 144, 0,
  1, 0, 144, 0,
  1, 0, 144, 0,
  1, 0, 176, 8192,
  0, 0, 160, 8192,
  0, 0, 160, 8192,
  0, 0, 160, 8192,
  0, 0, 160, 8192,
  1, 12, 3776, 8192,
  0, 0, 160, 8192,
  1, 0, 164, 8192,
  0, 0, 160, 8192,
  0, 0, 160, 8192,
  1, 0, 172, 8192,
  0, 0, 160, 8192,
  0, 0, 160, 8192,
  0, 0, 160, 8192,
  1, 0, 164, 8192,
  1, 0, 188, 8192,
  1, 0, 180, 8192,
  1, 0, 180, 8192,
  1, 0, 164, 8192,
  1, 0, 164, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 180, 8192,
  1, 0, 180, 8192,
  1, 0, 176, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 172, 8192,
  1, 0, 172, 8192,
  1, 0, 172, 8192,
  1, 0, 172, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 172, 8192,
  1, 0, 172, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 176, 8192,
  1, 0, 188, 8192,
  1, 0, 176, 8192,
  1, 0, 176, 8192,
  1, 0, 176, 8192,
  1, 0, 176, 8192,
  1, 0, 176, 8192,
  1, 0, 176, 8192,
  0, 0, 160, 8192,
  0, 0, 160, 8192,
  0, 0, 160, 8192,
  0, 0, 128, 8192,
  1, 0, 176, 8192,
  1, 0, 180, 8192,
  0, 0, 32, 4096,
  0, 0, 0, 4096,
  0, 0, 0, 4096,
  1, 0, 16, 4096,
  1, 0, 48, 4096,
  1, 0, 48, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 20, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 52, 4096,
  1, 0, 48, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  0, 0, 0, 4096,
  1, 0, 20, 4096,
  0, 0, 32, 4096,
  1, 0, 144, 0,
  0, 0, 128, 0,
  1, 0, 144, 0,
  1, 0, 144, 0,
  1, 0, 144, 0,
  1, 0, 144, 0,
  1, 0, 144, 0,
  1, 0, 144, 0,
  0, 0, 160, 8192,
  0, 0, 160, 8192,
  0, 0, 160, 8192,
  0, 0, 160, 8192,
  0, 0, 160, 8192,
  0, 0, 160, 8192,
  1, 0, 172, 8192,
  1, 0, 140, 8192,
  1, 0, 172, 8192,
  1, 0, 172, 8192,
  0, 0, 160, 8192,
  0, 0, 160, 8192,
  0, 0, 160, 8192,
  0, 0, 160, 8192,
  0, 0, 160, 8192,
  0, 0, 160, 8192,
  1, 0, 180, 8192,
  1, 0, 164, 8192,
  1, 0, 164, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 180, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 176, 8192,
  1, 0, 188, 8192,
  1, 0, 176, 8192,
  1, 0, 188, 8192,
  1, 0, 172, 8192,
  1, 0, 188, 8192,
  1, 0, 172, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 172, 8192,
  1, 0, 172, 8192,
  1, 0, 172, 8192,
  1, 0, 172, 8192,
  1, 0, 172, 8192,
  1, 0, 172, 8192,
  1, 0, 172, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 176, 8192,
  1, 0, 176, 8192,
  1, 0, 144, 8192,
  1, 0, 144, 8192,
  1, 0, 144, 8192,
  1, 0, 144, 8192,
  1, 0, 176, 8192,
  1, 0, 180, 8192,
  1, 0, 144, 8192,
  0, 0, 0, 4096,
  1, 0, 176, 8192,
  0, 0, 0, 4096,
  0, 0, 0, 4096,
  0, 0, 0, 4096,
  0, 0, 0, 4096,
  0, 0, 0, 4096,
  1, 0, 48, 4096,
  1, 0, 48, 4096,
  1, 0, 16, 4096,
  0, 0, 0, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 48, 4096,
  1, 0, 48, 4096,
  1, 0, 52, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 20, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 20, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  0, 0, 32, 4096,
  0, 0, 32, 4096,
  0, 0, 32, 4096,
  0, 0, 32, 4096,
  0, 0, 128, 0,
  0, 0, 128, 0,
  1, 0, 144, 0,
  1, 0, 144, 0,
  1, 0, 144, 0,
  1, 0, 144, 0,
  1, 0, 148, 0,
  0, 0, 160, 8192,
  0, 0, 160, 8192,
  0, 0, 160, 8192,
  0, 0, 160, 8192,
  0, 0, 160, 8192,
  1, 0, 172, 8192,
  0, 0, 128, 8192,
  0, 0, 128, 8192,
  1, 0, 172, 8192,
  0, 0, 160, 8192,
  0, 0, 160, 8192,
  0, 0, 160, 8192,
  0, 0, 160, 8192,
  0, 0, 160, 8192,
  0, 0, 160, 8192,
  1, 0, 164, 8192,
  0, 0, 160, 8192,
  1, 0, 164, 8192,
  1, 0, 180, 8192,
  1, 0, 180, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 176, 8192,
  1, 0, 188, 8192,
  1, 0, 180, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 180, 8192,
  1, 0, 188, 8192,
  1, 0, 180, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 172, 8192,
  1, 0, 172, 8192,
  1, 0, 172, 8192,
  1, 0, 172, 8192,
  1, 0, 172, 8192,
  1, 0, 172, 8192,
  1, 0, 172, 8192,
  1, 0, 188, 8192,
  1, 0, 176, 8192,
  1, 0, 176, 8192,
  1, 0, 176, 8192,
  1, 0, 176, 8192,
  1, 0, 176, 8192,
  1, 0, 144, 8192,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 144, 8192,
  0, 0, 0, 4096,
  0, 0, 0, 4096,
  0, 0, 0, 4096,
  0, 0, 0, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  0, 0, 0, 4096,
  0, 0, 0, 4096,
  1, 0, 48, 4096,
  0, 0, 32, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  0, 0, 0, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 48, 4096,
  1, 0, 48, 4096,
  1, 0, 16, 4096,
  1, 0, 28, 4096,
  1, 0, 20, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 48, 4096,
  1, 0, 48, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 48, 4096,
  1, 0, 48, 4096,
  0, 0, 32, 4096,
  0, 0, 32, 4096,
  0, 0, 32, 4096,
  0, 0, 128, 0,
  1, 0, 144, 0,
  1, 0, 144, 0,
  1, 0, 144, 0,
  1, 0, 144, 0,
  1, 0, 144, 0,
  1, 0, 156, 0 ;

 RAzi_angle =
  44.01, 44.82, 45.58, 46.3, 46.98, 47.63, 48.24, 48.83, 49.41, 49.96, 50.49, 
    50.99, 51.49, 51.98, 52.45, 52.9, 53.34, 53.78, 54.21, 54.62, 55.03, 
    55.42, 55.82, 56.21, 56.59, 56.95, 57.32, 57.68, 58.04, 58.4, 58.75, 
    59.09, 59.43, 59.78, 60.11, 60.44, 60.77, 61.1, 61.43, 61.74, 62.05, 
    62.35, 62.65, 62.92, 63.15, 63.3, 63.19, 61.14, -112.15, -113.72, 
    -113.78, -113.61, -113.35, -113.05, -112.73, -112.4, -112.05, -111.68, 
    -111.31, -110.94, -110.56, -110.16, -109.75, -109.34, -108.92, -108.49, 
    -108.05, -107.59, -107.12, -106.64, -106.15, -105.65, -105.12, -104.58, 
    -104.02, -103.45, -102.85, -102.22, -101.57, -100.9, -100.21, -99.48, 
    -98.71, -97.89, -97.06, -96.18, -95.23, -94.24, -93.18, -92.06, -90.87, 
    -89.58, -88.18, -86.68, -85.07, -83.32,
  43.76, 44.58, 45.34, 46.06, 46.73, 47.38, 48, 48.6, 49.17, 49.71, 50.25, 
    50.76, 51.27, 51.74, 52.21, 52.67, 53.12, 53.56, 53.98, 54.39, 54.8, 
    55.2, 55.6, 55.98, 56.36, 56.73, 57.11, 57.47, 57.83, 58.18, 58.53, 
    58.88, 59.23, 59.57, 59.9, 60.24, 60.58, 60.9, 61.22, 61.54, 61.85, 
    62.16, 62.46, 62.73, 62.96, 63.1, 62.98, 60.87, -112.23, -113.88, 
    -113.95, -113.77, -113.51, -113.21, -112.89, -112.55, -112.2, -111.84, 
    -111.47, -111.09, -110.7, -110.3, -109.89, -109.48, -109.06, -108.62, 
    -108.17, -107.71, -107.25, -106.76, -106.26, -105.74, -105.22, -104.68, 
    -104.12, -103.53, -102.92, -102.3, -101.66, -100.98, -100.27, -99.52, 
    -98.76, -97.95, -97.1, -96.2, -95.24, -94.25, -93.2, -92.06, -90.83, 
    -89.52, -88.14, -86.65, -85.01, -83.2,
  43.53, 44.34, 45.09, 45.81, 46.49, 47.14, 47.76, 48.35, 48.92, 49.48, 
    50.02, 50.53, 51.02, 51.5, 51.98, 52.44, 52.89, 53.32, 53.74, 54.16, 
    54.57, 54.97, 55.37, 55.75, 56.14, 56.52, 56.89, 57.25, 57.61, 57.97, 
    58.32, 58.67, 59.01, 59.35, 59.7, 60.04, 60.37, 60.69, 61.02, 61.34, 
    61.66, 61.96, 62.26, 62.53, 62.77, 62.91, 62.79, 60.75, -112.35, -114.05, 
    -114.11, -113.94, -113.68, -113.38, -113.05, -112.71, -112.36, -112, 
    -111.62, -111.24, -110.85, -110.45, -110.04, -109.62, -109.19, -108.75, 
    -108.3, -107.85, -107.37, -106.87, -106.37, -105.86, -105.34, -104.79, 
    -104.22, -103.63, -103.02, -102.39, -101.73, -101.04, -100.33, -99.6, 
    -98.82, -97.99, -97.12, -96.23, -95.28, -94.27, -93.19, -92.03, -90.81, 
    -89.51, -88.11, -86.58, -84.91, -83.11,
  43.27, 44.07, 44.84, 45.57, 46.24, 46.88, 47.5, 48.11, 48.68, 49.23, 49.76, 
    50.28, 50.78, 51.27, 51.74, 52.2, 52.64, 53.09, 53.52, 53.93, 54.34, 
    54.74, 55.14, 55.54, 55.92, 56.29, 56.66, 57.03, 57.4, 57.75, 58.1, 
    58.45, 58.8, 59.15, 59.49, 59.82, 60.16, 60.49, 60.82, 61.14, 61.45, 
    61.76, 62.06, 62.33, 62.56, 62.71, 62.58, 60.38, -112.55, -114.2, 
    -114.28, -114.1, -113.84, -113.54, -113.22, -112.88, -112.52, -112.15, 
    -111.77, -111.39, -111, -110.6, -110.18, -109.75, -109.33, -108.89, 
    -108.44, -107.97, -107.49, -107, -106.5, -105.98, -105.44, -104.88, 
    -104.32, -103.73, -103.11, -102.46, -101.8, -101.12, -100.41, -99.66, 
    -98.86, -98.03, -97.17, -96.27, -95.3, -94.27, -93.19, -92.04, -90.81, 
    -89.47, -88.04, -86.51, -84.86, -83.05,
  43.02, 43.84, 44.6, 45.31, 45.99, 46.64, 47.27, 47.86, 48.43, 48.98, 49.52, 
    50.04, 50.54, 51.02, 51.49, 51.96, 52.41, 52.85, 53.28, 53.69, 54.11, 
    54.52, 54.91, 55.3, 55.68, 56.06, 56.44, 56.81, 57.17, 57.53, 57.89, 
    58.24, 58.59, 58.93, 59.27, 59.61, 59.95, 60.29, 60.61, 60.93, 61.25, 
    61.57, 61.86, 62.13, 62.37, 62.52, 62.38, 60.19, -112.65, -114.38, 
    -114.46, -114.28, -114.02, -113.72, -113.39, -113.04, -112.68, -112.31, 
    -111.94, -111.55, -111.15, -110.74, -110.33, -109.91, -109.47, -109.02, 
    -108.56, -108.1, -107.62, -107.13, -106.61, -106.09, -105.55, -105, 
    -104.43, -103.82, -103.19, -102.56, -101.9, -101.2, -100.47, -99.71, 
    -98.92, -98.09, -97.21, -96.28, -95.3, -94.29, -93.21, -92.03, -90.77, 
    -89.43, -88.01, -86.48, -84.79, -82.92,
  42.78, 43.59, 44.34, 45.06, 45.74, 46.39, 47.01, 47.6, 48.18, 48.74, 49.28, 
    49.79, 50.29, 50.78, 51.26, 51.72, 52.17, 52.6, 53.04, 53.46, 53.88, 
    54.28, 54.67, 55.07, 55.46, 55.84, 56.21, 56.58, 56.95, 57.31, 57.67, 
    58.02, 58.36, 58.71, 59.06, 59.4, 59.74, 60.07, 60.4, 60.73, 61.05, 
    61.36, 61.66, 61.94, 62.18, 62.33, 62.2, 60.12, -112.91, -114.58, 
    -114.64, -114.47, -114.2, -113.9, -113.56, -113.21, -112.86, -112.49, 
    -112.1, -111.71, -111.31, -110.91, -110.49, -110.05, -109.61, -109.17, 
    -108.71, -108.24, -107.75, -107.25, -106.74, -106.22, -105.67, -105.1, 
    -104.52, -103.92, -103.3, -102.65, -101.97, -101.27, -100.54, -99.78, 
    -98.98, -98.13, -97.24, -96.33, -95.35, -94.31, -93.19, -92.01, -90.76, 
    -89.42, -87.97, -86.4, -84.69, -82.85,
  42.51, 43.32, 44.09, 44.81, 45.49, 46.13, 46.75, 47.36, 47.93, 48.49, 
    49.02, 49.54, 50.05, 50.54, 51.01, 51.47, 51.92, 52.37, 52.8, 53.22, 
    53.63, 54.04, 54.44, 54.84, 55.22, 55.6, 55.98, 56.36, 56.72, 57.08, 
    57.44, 57.79, 58.15, 58.5, 58.84, 59.18, 59.53, 59.87, 60.2, 60.52, 
    60.84, 61.16, 61.46, 61.74, 61.98, 62.13, 62.02, 59.86, -113.16, -114.78, 
    -114.84, -114.65, -114.38, -114.07, -113.74, -113.4, -113.03, -112.65, 
    -112.27, -111.88, -111.48, -111.06, -110.63, -110.2, -109.77, -109.32, 
    -108.85, -108.37, -107.88, -107.39, -106.87, -106.33, -105.78, -105.22, 
    -104.64, -104.03, -103.39, -102.73, -102.05, -101.36, -100.62, -99.84, 
    -99.03, -98.19, -97.3, -96.37, -95.36, -94.31, -93.2, -92.03, -90.76, 
    -89.38, -87.91, -86.35, -84.65, -82.77,
  42.26, 43.08, 43.84, 44.55, 45.23, 45.88, 46.51, 47.1, 47.67, 48.23, 48.77, 
    49.3, 49.8, 50.28, 50.76, 51.23, 51.68, 52.12, 52.55, 52.97, 53.39, 
    53.81, 54.21, 54.6, 54.99, 55.37, 55.75, 56.12, 56.49, 56.85, 57.22, 
    57.58, 57.93, 58.27, 58.62, 58.97, 59.32, 59.65, 59.98, 60.31, 60.64, 
    60.96, 61.26, 61.54, 61.79, 61.95, 61.84, 59.77, -113.3, -114.99, 
    -115.04, -114.85, -114.58, -114.27, -113.93, -113.57, -113.2, -112.83, 
    -112.45, -112.05, -111.64, -111.22, -110.8, -110.37, -109.92, -109.46, 
    -108.99, -108.52, -108.03, -107.52, -106.99, -106.45, -105.91, -105.34, 
    -104.74, -104.13, -103.49, -102.84, -102.15, -101.44, -100.68, -99.91, 
    -99.1, -98.25, -97.34, -96.39, -95.4, -94.35, -93.22, -92, -90.71, 
    -89.34, -87.89, -86.31, -84.56, -82.65,
  42.01, 42.81, 43.57, 44.29, 44.98, 45.63, 46.24, 46.84, 47.42, 47.99, 
    48.52, 49.03, 49.54, 50.03, 50.52, 50.98, 51.43, 51.87, 52.31, 52.74, 
    53.15, 53.56, 53.96, 54.36, 54.75, 55.14, 55.51, 55.89, 56.26, 56.63, 
    56.99, 57.34, 57.7, 58.05, 58.41, 58.75, 59.09, 59.43, 59.77, 60.11, 
    60.43, 60.75, 61.05, 61.34, 61.59, 61.75, 61.66, 59.65, -113.63, -115.2, 
    -115.24, -115.05, -114.77, -114.45, -114.11, -113.76, -113.39, -113.01, 
    -112.61, -112.21, -111.81, -111.39, -110.96, -110.52, -110.07, -109.61, 
    -109.15, -108.66, -108.16, -107.65, -107.13, -106.59, -106.03, -105.45, 
    -104.85, -104.24, -103.6, -102.93, -102.23, -101.51, -100.77, -99.99, 
    -99.16, -98.29, -97.37, -96.43, -95.43, -94.36, -93.21, -92, -90.71, 
    -89.33, -87.84, -86.22, -84.47, -82.59,
  41.73, 42.55, 43.31, 44.03, 44.71, 45.36, 45.98, 46.59, 47.16, 47.72, 
    48.25, 48.78, 49.29, 49.78, 50.26, 50.72, 51.18, 51.63, 52.06, 52.48, 
    52.9, 53.31, 53.72, 54.12, 54.51, 54.89, 55.27, 55.66, 56.03, 56.39, 
    56.75, 57.12, 57.47, 57.82, 58.17, 58.52, 58.87, 59.22, 59.55, 59.88, 
    60.21, 60.53, 60.84, 61.13, 61.38, 61.54, 61.43, 59.3, -113.76, -115.38, 
    -115.42, -115.23, -114.95, -114.64, -114.3, -113.94, -113.56, -113.18, 
    -112.79, -112.39, -111.98, -111.55, -111.12, -110.68, -110.23, -109.76, 
    -109.28, -108.8, -108.3, -107.79, -107.26, -106.71, -106.14, -105.57, 
    -104.97, -104.34, -103.69, -103.01, -102.32, -101.61, -100.85, -100.05, 
    -99.21, -98.35, -97.44, -96.47, -95.44, -94.36, -93.22, -92.01, -90.69, 
    -89.27, -87.77, -86.17, -84.42, -82.49,
  41.49, 42.3, 43.05, 43.76, 44.45, 45.11, 45.73, 46.33, 46.9, 47.46, 48.01, 
    48.53, 49.03, 49.52, 50, 50.47, 50.93, 51.37, 51.8, 52.23, 52.66, 53.07, 
    53.47, 53.87, 54.26, 54.66, 55.04, 55.41, 55.78, 56.16, 56.52, 56.88, 
    57.24, 57.59, 57.95, 58.3, 58.65, 58.99, 59.33, 59.66, 60, 60.32, 60.63, 
    60.92, 61.17, 61.34, 61.24, 59.25, -113.96, -115.59, -115.63, -115.43, 
    -115.16, -114.83, -114.49, -114.12, -113.75, -113.37, -112.97, -112.56, 
    -112.14, -111.72, -111.29, -110.84, -110.38, -109.91, -109.44, -108.95, 
    -108.45, -107.92, -107.38, -106.84, -106.28, -105.69, -105.08, -104.45, 
    -103.8, -103.13, -102.42, -101.68, -100.91, -100.12, -99.29, -98.4, 
    -97.47, -96.5, -95.48, -94.4, -93.23, -91.98, -90.66, -89.25, -87.75, 
    -86.1, -84.31, -82.36,
  41.21, 42.01, 42.77, 43.5, 44.19, 44.83, 45.45, 46.06, 46.64, 47.2, 47.74, 
    48.25, 48.76, 49.26, 49.75, 50.21, 50.67, 51.11, 51.56, 51.99, 52.4, 
    52.81, 53.22, 53.63, 54.02, 54.41, 54.79, 55.17, 55.55, 55.92, 56.28, 
    56.64, 57, 57.36, 57.72, 58.07, 58.42, 58.76, 59.11, 59.44, 59.77, 60.1, 
    60.41, 60.71, 60.96, 61.13, 61.04, 59.06, -114.26, -115.8, -115.83, 
    -115.64, -115.35, -115.02, -114.68, -114.32, -113.94, -113.54, -113.14, 
    -112.74, -112.32, -111.9, -111.45, -111, -110.54, -110.08, -109.6, 
    -109.1, -108.58, -108.06, -107.53, -106.98, -106.4, -105.8, -105.2, 
    -104.57, -103.91, -103.22, -102.5, -101.77, -101, -100.2, -99.34, -98.45, 
    -97.52, -96.55, -95.51, -94.4, -93.22, -91.98, -90.66, -89.23, -87.68, 
    -86.02, -84.24, -82.3 ;

 RFlag =
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888 ;

 RR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 12, 11, 9, 10, 7, 8, 0, 0, 0, 0, 6, 5, 7, 
    8, 6, 6, 5, 6, 8, 9, 8, 9, 13, 12, 11, 8, 6, 8, 7, 6, 0, 0, 0, 0, 0, 0, 
    0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 0, 0, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 12, 16, 10, 6, 11, 10, 6, 6, 5, 6, 6, 9, 10, 
    12, 7, 8, 6, 7, 6, 7, 7, 7, 7, 7, 6, 10, 10, 12, 9, 7, 5, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 4, 13, 12, 11, 7, 11, 7, 14, 8, 6, 7, 5, 6, 6, 6, 
    6, 8, 10, 8, 7, 6, 0, 0, 0, 5, 7, 6, 6, 8, 7, 8, 8, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 7, 6, 15, 9, 5, 8, 7, 6, 7, 8, 9, 8, 6, 6, 9, 7, 9, 9, 
    7, 5, 10, 0, 0, 5, 7, 0, 8, 8, 7, 5, 5, 6, 6, 5, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 9, 14, 7, 5, 11, 0, 0, 9, 8, 8, 6, 6, 7, 12, 26, 
    12, 7, 11, 9, 7, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, 0, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 5, 11, 6, 8, 25, 13, 8, 6, 6, 7, 6, 5, 6, 6, 12, 20, 
    7, 0, 7, 6, 8, 0, 0, 0, 0, 0, 0, 0, 5, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 6, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 9, 7, 9, 7, 5, 14, 12, 5, 5, 7, 8, 6, 5, 14, 19, 15, 6, 
    9, 7, 6, 0, 0, 0, 0, 0, 0, 6, 7, 7, 6, 0, 0, 5, 5, 0, 0, 9, 15, 12, 11, 
    8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0, 0, 0, 0, 0, 10, 5, 8, 5, 6, 8, 7, 5, 0, 0, 0, 0, 0, 6, 14, 11, 8, 6, 7, 
    6, 0, 6, 5, 0, 0, 0, 0, 0, 7, 7, 6, 7, 0, 0, 5, 0, 17, 20, 18, 14, 11, 
    11, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0, 0, 0, 0, 6, 6, 5, 14, 5, 0, 0, 0, 5, 0, 0, 0, 7, 6, 8, 23, 9, 7, 5, 6, 
    7, 0, 19, 6, 0, 0, 0, 0, 0, 6, 9, 8, 21, 17, 6, 14, 20, 15, 5, 5, 6, 5, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0, 0, 0, 6, 17, 6, 7, 0, 0, 0, 0, 5, 5, 0, 0, 0, 5, 0, 0, 5, 5, 0, 7, 6, 0, 
    0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 6, 0, 6, 9, 0, 8, 6, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 10, 19, 5, 0, 0, 0, 0, 0, 5, 6, 0, 0, 0, 5, 0, 5, 6, 6, 8, 0, 0, 
    7, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, _, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 7, 5, 0, 2, 3, 0, 0, 0, 5, 0, 0, 0, 0, 6, 0, 0, 7, 5, 8, 0, 7, 9, 
    0, 0, 6, 7, 6, 0, 0, 0, 0, 7, 8, 5, 0, 6, 8, 9, 7, 0, 0, 0, 0, 0, 0, _, 
    _, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 RWP =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 13, 7, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    7, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 0, 0, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 10, 10, 11, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 8, 14, 17, 13, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 13, 10, 12, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 15, 13, 13, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, 0, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 10, 17, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 12, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 11, 11, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 10, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, _, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 3, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, 
    _, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 SFR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 0, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 0, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 SIce =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, 38, 24, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 40, 56, 66, 78, 78, 78, _, _, 82, 78, 68, 
    60, 60,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, 0, 0, 0, 0, 0, 0, 0, 50, 0, 50, 0, 52, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 40, 56, 66, 76, 80, 76, 78, 80, 84, 80, 
    74, 66, 64,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, 0, 0, 0, 0, 0, 0, 0, 0, 54, 56, 58, 
    56, 0, 0, 42, 0, 0, 0, 0, 0, 0, 0, 42, 58, 72, 76, 76, 80, 82, 82, 84, 
    78, 78, 74, 68,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, 0, 0, 0, 0, 0, 0, 0, 58, 60, 62, 0, 
    0, 0, 0, 48, 0, 0, 0, 0, 0, 0, 0, 46, 58, 70, 76, 78, 78, 78, 80, 82, 82, 
    80, 78, 74,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, 0, _, 0, 0, 0, 0, 62, 0, 0, 62, 0, 0, 
    56, 0, 50, 0, 0, 0, 0, 0, 26, 40, 56, 60, 68, 78, 78, 78, 82, 82, 84, 84, 
    82, 76, 76,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, 0, 0, 0, 0, 0, 0, 0, 64, 62, 62, 62, 58, 
    0, 0, 52, 52, 0, 0, 0, 36, 0, 42, 52, 64, 62, 68, 76, 78, 82, 82, 84, 88, 
    88, 88, 82, 80,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, 0, 48, 0, 0, 58, 64, 66, 66, 62, 62, 60, 
    56, 52, 50, 50, 52, 50, 50, 48, 48, 46, 56, 56, 58, 64, 72, 76, 80, 82, 
    84, 84, 88, 90, 92, 84, 84,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, 0, 0, 0, 56, 0, 66, 68, 68, 64, 62, 0, 
    52, 48, 46, 48, 52, 54, 54, 54, 54, 54, 56, 60, 62, 68, 70, 76, 78, 82, 
    84, 88, 90, 94, 92, 88, 84,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, 0, 0, 0, 0, 0, 0, 0, 66, 0, 70, 70, 64, 0, 0, 52, 
    48, 46, 48, 52, 56, 60, 60, 62, 62, 62, 62, 66, 68, 68, 74, 76, 80, 86, 
    88, 90, 94, 90, 86, 82,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, 0, 0, 0, 0, 0, 0, 64, 68, 70, 72, 70, 66, 64, 58, 
    54, 48, 46, 48, 52, 58, 62, 64, 64, 66, 66, 66, 68, 68, 68, 74, 78, 82, 
    84, 86, 92, 90, 90, 88, 84,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, 0, _, 60, 0, 0, 0, 0, 0, 0, 64, 68, 70, 72, 72, 72, 68, 64, 
    60, 52, 48, 46, 50, 56, 62, 66, 66, 68, 68, 68, 66, 68, 68, 68, 74, 78, 
    82, 84, 88, 92, 90, 94, 90, 88,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 70, 
    72, _, 72, 0, 0, 54, 0, 0, 0, 0, 0, 60, 64, 68, 70, 72, 72, 72, 72, 68, 
    62, 56, 50, 44, 46, 52, 58, 64, 68, 68, 70, 68, 68, 68, 68, 70, 70, 74, 
    78, 82, 84, 90, 96, 94, 96, 92, 88 ;

 SIce_FY =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, 38, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 40, 56, 66, 78, 78, 78, _, _, 82, 78, 68, 
    60, 60,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, 0, 0, 0, 0, 0, 0, 0, 50, 0, 50, 0, 52, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 40, 56, 66, 76, 80, 76, 78, 80, 84, 80, 
    74, 66, 64,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, 0, 0, 0, 0, 0, 0, 0, 0, 54, 56, 58, 
    56, 0, 0, 42, 0, 0, 0, 0, 0, 0, 0, 42, 58, 72, 76, 76, 80, 82, 82, 84, 
    78, 78, 74, 68,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, 0, 0, 0, 0, 0, 0, 0, 58, 60, 62, 0, 
    0, 0, 0, 48, 0, 0, 0, 0, 0, 0, 0, 46, 58, 70, 76, 78, 78, 78, 80, 82, 82, 
    80, 78, 74,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, 0, _, 0, 0, 0, 0, 62, 0, 0, 62, 0, 0, 
    56, 0, 50, 0, 0, 0, 0, 0, 0, 40, 56, 60, 68, 78, 78, 78, 82, 82, 84, 84, 
    82, 76, 76,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, 0, 0, 0, 0, 0, 0, 0, 64, 62, 62, 62, 58, 
    0, 0, 52, 52, 0, 0, 0, 36, 0, 42, 52, 64, 62, 68, 76, 78, 82, 82, 84, 88, 
    88, 88, 82, 80,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, 0, 48, 0, 0, 58, 64, 66, 66, 62, 62, 60, 
    56, 52, 50, 50, 52, 50, 50, 48, 48, 46, 56, 56, 58, 64, 72, 76, 80, 82, 
    84, 84, 88, 90, 92, 84, 84,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, 0, 0, 0, 56, 0, 66, 68, 68, 64, 62, 0, 
    52, 48, 46, 48, 52, 54, 54, 54, 54, 54, 56, 60, 62, 68, 70, 76, 78, 82, 
    84, 88, 90, 94, 92, 88, 84,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, 0, 0, 0, 0, 0, 0, 0, 66, 0, 70, 70, 64, 0, 0, 52, 
    48, 46, 48, 52, 56, 60, 60, 62, 62, 62, 62, 66, 68, 68, 74, 76, 80, 86, 
    88, 90, 94, 90, 86, 82,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, 0, 0, 0, 0, 0, 0, 64, 68, 70, 72, 70, 66, 64, 58, 
    54, 48, 46, 48, 52, 58, 62, 64, 64, 66, 66, 66, 68, 68, 68, 74, 78, 82, 
    84, 86, 92, 90, 90, 88, 84,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, 0, _, 60, 0, 0, 0, 0, 0, 0, 64, 68, 70, 72, 72, 72, 68, 64, 
    60, 52, 48, 46, 50, 56, 62, 66, 66, 68, 68, 68, 66, 68, 68, 68, 74, 78, 
    82, 84, 88, 92, 90, 94, 90, 88,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 70, 
    72, _, 72, 0, 0, 54, 0, 0, 0, 0, 0, 60, 64, 68, 70, 72, 72, 72, 72, 68, 
    62, 56, 50, 44, 46, 52, 58, 64, 68, 68, 70, 68, 68, 68, 68, 70, 70, 74, 
    78, 82, 84, 90, 96, 94, 96, 92, 88 ;

 SIce_MY =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, 0, 0, 0, 0, 0,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, 0, _, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 25, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, 0, _, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 0, 
    0, _, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SWE =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 0, 0, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, 0, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, _, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, 
    _, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 SWP =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 SZ_angle =
  43.11, 43.21, 43.31, 43.41, 43.51, 43.6, 43.68, 43.77, 43.85, 43.93, 44.01, 
    44.08, 44.15, 44.23, 44.3, 44.36, 44.43, 44.5, 44.56, 44.62, 44.68, 
    44.74, 44.8, 44.86, 44.92, 44.98, 45.03, 45.09, 45.14, 45.2, 45.25, 45.3, 
    45.36, 45.41, 45.46, 45.51, 45.57, 45.62, 45.67, 45.72, 45.77, 45.82, 
    45.87, 45.93, 45.98, 46.03, 46.08, 46.13, 46.19, 46.24, 46.29, 46.35, 
    46.4, 46.46, 46.51, 46.57, 46.62, 46.68, 46.74, 46.8, 46.86, 46.92, 
    46.98, 47.05, 47.11, 47.18, 47.24, 47.31, 47.39, 47.46, 47.53, 47.61, 
    47.69, 47.77, 47.86, 47.94, 48.04, 48.13, 48.23, 48.33, 48.44, 48.55, 
    48.67, 48.79, 48.92, 49.06, 49.2, 49.36, 49.52, 49.7, 49.89, 50.1, 50.32, 
    50.57, 50.84, 51.13,
  43.26, 43.37, 43.47, 43.56, 43.66, 43.75, 43.83, 43.92, 44, 44.08, 44.16, 
    44.23, 44.31, 44.38, 44.45, 44.52, 44.58, 44.65, 44.71, 44.77, 44.83, 
    44.9, 44.96, 45.01, 45.07, 45.13, 45.18, 45.24, 45.29, 45.35, 45.4, 
    45.45, 45.51, 45.56, 45.61, 45.66, 45.72, 45.77, 45.82, 45.87, 45.92, 
    45.97, 46.02, 46.07, 46.12, 46.18, 46.23, 46.28, 46.33, 46.39, 46.44, 
    46.49, 46.55, 46.6, 46.66, 46.71, 46.77, 46.83, 46.89, 46.94, 47, 47.07, 
    47.13, 47.19, 47.26, 47.32, 47.39, 47.46, 47.53, 47.6, 47.68, 47.76, 
    47.83, 47.91, 48, 48.09, 48.18, 48.27, 48.37, 48.47, 48.58, 48.69, 48.81, 
    48.93, 49.06, 49.2, 49.34, 49.5, 49.66, 49.84, 50.03, 50.24, 50.46, 50.7, 
    50.97, 51.27,
  43.41, 43.52, 43.62, 43.71, 43.81, 43.9, 43.99, 44.07, 44.15, 44.23, 44.31, 
    44.39, 44.46, 44.53, 44.6, 44.67, 44.73, 44.8, 44.86, 44.92, 44.98, 
    45.04, 45.1, 45.16, 45.22, 45.28, 45.33, 45.39, 45.44, 45.5, 45.55, 45.6, 
    45.66, 45.71, 45.76, 45.81, 45.86, 45.91, 45.97, 46.02, 46.07, 46.12, 
    46.17, 46.22, 46.27, 46.32, 46.38, 46.43, 46.48, 46.53, 46.59, 46.64, 
    46.69, 46.75, 46.8, 46.86, 46.92, 46.97, 47.03, 47.09, 47.15, 47.21, 
    47.27, 47.34, 47.4, 47.47, 47.53, 47.6, 47.67, 47.75, 47.82, 47.9, 47.98, 
    48.06, 48.14, 48.23, 48.32, 48.41, 48.51, 48.61, 48.72, 48.83, 48.95, 
    49.07, 49.2, 49.34, 49.48, 49.63, 49.8, 49.98, 50.17, 50.37, 50.59, 
    50.84, 51.11, 51.41,
  43.56, 43.67, 43.77, 43.87, 43.96, 44.05, 44.14, 44.22, 44.3, 44.38, 44.46, 
    44.54, 44.61, 44.68, 44.75, 44.82, 44.88, 44.95, 45.01, 45.07, 45.13, 
    45.19, 45.25, 45.31, 45.37, 45.43, 45.48, 45.54, 45.59, 45.65, 45.7, 
    45.75, 45.8, 45.86, 45.91, 45.96, 46.01, 46.06, 46.11, 46.17, 46.22, 
    46.27, 46.32, 46.37, 46.42, 46.47, 46.52, 46.57, 46.63, 46.68, 46.73, 
    46.79, 46.84, 46.9, 46.95, 47, 47.06, 47.12, 47.18, 47.24, 47.29, 47.36, 
    47.42, 47.48, 47.55, 47.61, 47.68, 47.75, 47.82, 47.89, 47.96, 48.04, 
    48.12, 48.2, 48.28, 48.37, 48.46, 48.56, 48.66, 48.76, 48.86, 48.97, 
    49.09, 49.21, 49.34, 49.47, 49.62, 49.77, 49.94, 50.11, 50.3, 50.51, 
    50.73, 50.97, 51.24, 51.53,
  43.72, 43.82, 43.92, 44.02, 44.11, 44.2, 44.29, 44.37, 44.46, 44.53, 44.61, 
    44.69, 44.76, 44.83, 44.9, 44.97, 45.03, 45.1, 45.16, 45.22, 45.28, 
    45.35, 45.4, 45.46, 45.52, 45.58, 45.63, 45.69, 45.74, 45.79, 45.85, 
    45.9, 45.95, 46.01, 46.06, 46.11, 46.16, 46.21, 46.26, 46.31, 46.36, 
    46.42, 46.47, 46.52, 46.57, 46.62, 46.67, 46.72, 46.77, 46.83, 46.88, 
    46.93, 46.99, 47.04, 47.1, 47.15, 47.21, 47.26, 47.32, 47.38, 47.44, 
    47.5, 47.56, 47.63, 47.69, 47.76, 47.82, 47.89, 47.96, 48.03, 48.11, 
    48.19, 48.26, 48.34, 48.43, 48.52, 48.61, 48.7, 48.8, 48.9, 49, 49.11, 
    49.23, 49.35, 49.48, 49.62, 49.76, 49.91, 50.07, 50.25, 50.44, 50.65, 
    50.87, 51.11, 51.37, 51.68,
  43.87, 43.97, 44.07, 44.17, 44.26, 44.35, 44.44, 44.52, 44.61, 44.69, 
    44.76, 44.84, 44.91, 44.98, 45.05, 45.12, 45.19, 45.25, 45.31, 45.38, 
    45.44, 45.5, 45.55, 45.61, 45.67, 45.73, 45.78, 45.84, 45.89, 45.94, 46, 
    46.05, 46.1, 46.15, 46.21, 46.26, 46.31, 46.36, 46.41, 46.46, 46.51, 
    46.56, 46.61, 46.66, 46.72, 46.77, 46.82, 46.87, 46.92, 46.97, 47.03, 
    47.08, 47.13, 47.19, 47.24, 47.3, 47.35, 47.41, 47.47, 47.53, 47.59, 
    47.65, 47.71, 47.77, 47.84, 47.9, 47.97, 48.04, 48.11, 48.18, 48.25, 
    48.33, 48.41, 48.49, 48.57, 48.66, 48.75, 48.84, 48.94, 49.04, 49.14, 
    49.25, 49.37, 49.49, 49.62, 49.76, 49.9, 50.05, 50.22, 50.39, 50.58, 
    50.78, 51, 51.24, 51.51, 51.81,
  44.02, 44.12, 44.23, 44.32, 44.42, 44.51, 44.59, 44.68, 44.76, 44.84, 
    44.91, 44.99, 45.06, 45.13, 45.2, 45.27, 45.34, 45.4, 45.46, 45.53, 
    45.59, 45.65, 45.7, 45.76, 45.82, 45.88, 45.93, 45.99, 46.04, 46.09, 
    46.15, 46.2, 46.25, 46.3, 46.35, 46.41, 46.46, 46.51, 46.56, 46.61, 
    46.66, 46.71, 46.76, 46.81, 46.86, 46.91, 46.96, 47.02, 47.07, 47.12, 
    47.17, 47.23, 47.28, 47.33, 47.39, 47.44, 47.5, 47.56, 47.61, 47.67, 
    47.73, 47.79, 47.85, 47.92, 47.98, 48.04, 48.11, 48.18, 48.25, 48.32, 
    48.4, 48.47, 48.55, 48.63, 48.71, 48.8, 48.89, 48.98, 49.08, 49.18, 
    49.28, 49.4, 49.51, 49.63, 49.76, 49.89, 50.04, 50.19, 50.35, 50.53, 
    50.71, 50.92, 51.14, 51.38, 51.64, 51.94,
  44.17, 44.28, 44.38, 44.47, 44.57, 44.66, 44.75, 44.83, 44.91, 44.99, 
    45.07, 45.14, 45.21, 45.28, 45.35, 45.42, 45.49, 45.55, 45.61, 45.67, 
    45.74, 45.8, 45.86, 45.91, 45.97, 46.03, 46.08, 46.14, 46.19, 46.24, 
    46.3, 46.35, 46.4, 46.45, 46.5, 46.56, 46.61, 46.66, 46.71, 46.76, 46.81, 
    46.86, 46.91, 46.96, 47.01, 47.06, 47.11, 47.16, 47.21, 47.27, 47.32, 
    47.37, 47.43, 47.48, 47.54, 47.59, 47.65, 47.7, 47.76, 47.82, 47.88, 
    47.94, 48, 48.06, 48.13, 48.19, 48.26, 48.32, 48.39, 48.47, 48.54, 48.62, 
    48.69, 48.77, 48.86, 48.94, 49.03, 49.13, 49.22, 49.32, 49.43, 49.54, 
    49.65, 49.77, 49.9, 50.04, 50.18, 50.33, 50.49, 50.67, 50.86, 51.06, 
    51.27, 51.51, 51.78, 52.08,
  44.33, 44.43, 44.53, 44.63, 44.72, 44.81, 44.9, 44.98, 45.06, 45.14, 45.22, 
    45.29, 45.36, 45.44, 45.51, 45.57, 45.64, 45.7, 45.76, 45.83, 45.89, 
    45.95, 46, 46.06, 46.12, 46.18, 46.23, 46.28, 46.34, 46.39, 46.45, 46.5, 
    46.55, 46.6, 46.65, 46.7, 46.75, 46.81, 46.86, 46.91, 46.96, 47.01, 
    47.06, 47.11, 47.16, 47.21, 47.26, 47.31, 47.36, 47.42, 47.47, 47.52, 
    47.57, 47.63, 47.68, 47.74, 47.79, 47.85, 47.91, 47.96, 48.02, 48.08, 
    48.14, 48.21, 48.27, 48.34, 48.4, 48.47, 48.54, 48.61, 48.68, 48.76, 
    48.84, 48.92, 49, 49.09, 49.17, 49.27, 49.37, 49.47, 49.57, 49.68, 49.79, 
    49.92, 50.04, 50.18, 50.32, 50.47, 50.63, 50.81, 50.99, 51.19, 51.41, 
    51.65, 51.92, 52.21,
  44.48, 44.58, 44.68, 44.78, 44.87, 44.96, 45.05, 45.13, 45.21, 45.29, 
    45.37, 45.44, 45.52, 45.59, 45.66, 45.72, 45.79, 45.85, 45.92, 45.98, 
    46.04, 46.1, 46.16, 46.21, 46.27, 46.32, 46.38, 46.44, 46.49, 46.54, 
    46.59, 46.65, 46.7, 46.75, 46.8, 46.85, 46.9, 46.95, 47, 47.05, 47.1, 
    47.16, 47.21, 47.26, 47.31, 47.36, 47.41, 47.46, 47.51, 47.56, 47.61, 
    47.67, 47.72, 47.77, 47.83, 47.88, 47.94, 48, 48.05, 48.11, 48.17, 48.23, 
    48.29, 48.35, 48.41, 48.48, 48.55, 48.61, 48.68, 48.75, 48.83, 48.9, 
    48.98, 49.06, 49.14, 49.23, 49.32, 49.41, 49.51, 49.61, 49.71, 49.82, 
    49.94, 50.05, 50.18, 50.32, 50.46, 50.61, 50.77, 50.94, 51.13, 51.33, 
    51.55, 51.79, 52.05, 52.34,
  44.63, 44.73, 44.83, 44.93, 45.02, 45.11, 45.2, 45.28, 45.36, 45.44, 45.52, 
    45.6, 45.67, 45.74, 45.81, 45.87, 45.94, 46, 46.06, 46.13, 46.19, 46.25, 
    46.31, 46.36, 46.42, 46.48, 46.53, 46.58, 46.64, 46.69, 46.74, 46.8, 
    46.85, 46.9, 46.95, 47, 47.05, 47.1, 47.15, 47.2, 47.25, 47.3, 47.35, 
    47.4, 47.45, 47.5, 47.56, 47.61, 47.66, 47.71, 47.76, 47.81, 47.87, 
    47.92, 47.98, 48.03, 48.09, 48.14, 48.2, 48.26, 48.32, 48.37, 48.43, 
    48.5, 48.56, 48.63, 48.69, 48.76, 48.83, 48.9, 48.97, 49.05, 49.12, 49.2, 
    49.29, 49.37, 49.46, 49.55, 49.65, 49.75, 49.85, 49.96, 50.08, 50.2, 
    50.32, 50.46, 50.6, 50.75, 50.91, 51.08, 51.27, 51.47, 51.68, 51.92, 
    52.19, 52.48,
  44.78, 44.88, 44.98, 45.08, 45.18, 45.27, 45.35, 45.44, 45.52, 45.6, 45.67, 
    45.75, 45.82, 45.89, 45.96, 46.02, 46.09, 46.15, 46.22, 46.28, 46.34, 
    46.4, 46.46, 46.51, 46.57, 46.62, 46.68, 46.73, 46.79, 46.84, 46.89, 
    46.95, 47, 47.05, 47.1, 47.15, 47.2, 47.25, 47.3, 47.35, 47.4, 47.45, 
    47.5, 47.55, 47.6, 47.65, 47.7, 47.75, 47.81, 47.86, 47.91, 47.96, 48.01, 
    48.07, 48.12, 48.18, 48.23, 48.29, 48.35, 48.4, 48.46, 48.52, 48.58, 
    48.64, 48.71, 48.77, 48.84, 48.9, 48.97, 49.04, 49.12, 49.19, 49.27, 
    49.35, 49.43, 49.52, 49.6, 49.7, 49.79, 49.89, 49.99, 50.1, 50.22, 50.34, 
    50.46, 50.59, 50.74, 50.89, 51.05, 51.22, 51.4, 51.61, 51.82, 52.06, 
    52.32, 52.61 ;

 ScanTime_UTC = 5258.00048828125, 5261.00048828125, 5264.00048828125, 
    5266.00048828125, 5269.00048828125, 5272.00048828125, 5274.00048828125, 
    5277.00048828125, 5280.00048828125, 5282.00048828125, 5285.00048828125, 
    5288.00048828125 ;

 ScanTime_dom = 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30 ;

 ScanTime_doy = 181, 181, 181, 181, 181, 181, 181, 181, 181, 181, 181, 181 ;

 ScanTime_hour = 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1 ;

 ScanTime_minute = 27, 27, 27, 27, 27, 27, 27, 27, 28, 28, 28, 28 ;

 ScanTime_month = 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6 ;

 ScanTime_second = 38, 41, 44, 46, 49, 52, 54, 57, 0, 2, 5, 8 ;

 ScanTime_year = 2021, 2021, 2021, 2021, 2021, 2021, 2021, 2021, 2021, 2021, 
    2021, 2021 ;

 Sfc_type =
  2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 2, 2, 1, 1, 1, 1, 1,
  2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 0, 1, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 
    0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 0, 0, 
    0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 0, 2, 0, 0, 0, 0, 1, 0, 0, 1, 0, 0, 
    1, 0, 1, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 0, 
    0, 1, 1, 0, 0, 0, 1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 0, 1, 0, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 0, 0, 0, 1, 0, 1, 1, 1, 1, 1, 0, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 0, 0, 0, 0, 0, 0, 0, 1, 0, 1, 1, 1, 0, 0, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 0, 2, 1, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 1, 
    1, 2, 1, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1 ;

 Snow =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 0, 0, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, 0, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, _, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, 
    _, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 SnowGS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 0, 0, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, 0, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, _, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, 
    _, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 SurfM =
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888 ;

 SurfP =
  9796, 9796, 9832, 9327, 9120, 9072, 8772, 8811, 8788, 8858, 8491, 8333, 
    8423, 8729, 8765, 9409, 9591, 8966, 8772, 8620, 9241, 9769, 10004, 10018, 
    9997, 9980, 9616, 9577, 9681, 9877, 9844, 9990, 10018, 10018, 10018, 
    10018, 10018, 10018, 10018, 10018, 10018, 10018, 10018, 10018, 10018, 
    10018, 10018, 10018, 10018, 10018, 10018, 10018, 10018, 10018, 10018, 
    10018, 10018, 10018, 10046, 9930, 9930, 10084, 10084, 10084, 10084, 
    10084, 10084, 10084, 10084, 10084, 10084, 10084, 10084, 10084, 10084, 
    10084, 10084, 10084, 10084, 10084, 10084, 10084, 10084, 10084, 10084, 
    10084, 9930, 9930, 10084, 10027, 9976, 9930, 9930, 9930, 9930, 9930,
  9796, 9824, 9784, 9280, 9310, 8952, 8893, 8802, 8736, 8765, 8585, 8419, 
    8371, 8683, 8750, 9699, 9783, 9135, 8682, 8699, 9443, 9924, 10007, 10018, 
    10018, 9987, 9897, 9587, 9776, 9870, 9952, 10015, 10018, 10018, 10018, 
    10018, 10018, 10018, 10018, 10018, 10018, 10018, 10018, 10018, 10018, 
    10018, 10018, 10018, 10018, 10018, 10018, 10018, 10018, 10018, 10018, 
    10018, 10018, 10018, 10046, 10097, 10084, 10084, 10084, 10084, 10084, 
    10084, 10084, 10084, 10084, 10084, 10084, 10084, 10084, 10084, 10084, 
    10084, 10084, 10084, 10084, 10084, 10084, 10084, 10084, 10084, 10084, 
    10084, 10084, 9930, 10084, 10084, 9930, 9930, 9930, 9930, 9930, 9930,
  9796, 9824, 9574, 9156, 9014, 9027, 8869, 8801, 8770, 8765, 8452, 8450, 
    8471, 8609, 9177, 9546, 9762, 9458, 8812, 8805, 9724, 9999, 10002, 10018, 
    10018, 10018, 9980, 9794, 9811, 9918, 9990, 9983, 9969, 10018, 10018, 
    10018, 10018, 10018, 10018, 10018, 10018, 10018, 10018, 10018, 10018, 
    10018, 10018, 10018, 10018, 10018, 10018, 10018, 10018, 10018, 10018, 
    10046, 10046, 10046, 10054, 10084, 10130, 10084, 10084, 10084, 10084, 
    10084, 10084, 10084, 10084, 10084, 10084, 10084, 10084, 10084, 10084, 
    10084, 10084, 10084, 10084, 10084, 10084, 10084, 10084, 10084, 10084, 
    10084, 10084, 10084, 9930, 10084, 9930, 9930, 9930, 9930, 9930, 9930,
  9796, 9832, 9671, 8824, 8956, 8781, 8838, 8745, 8906, 8600, 8391, 8598, 
    8662, 8609, 9143, 9421, 9553, 9592, 8750, 9393, 9906, 9992, 10018, 10018, 
    10018, 10018, 10010, 9987, 9946, 9835, 10008, 9976, 10008, 10014, 10018, 
    10018, 10018, 10018, 10018, 10018, 10018, 10018, 10018, 10018, 10018, 
    10018, 10018, 9976, 10018, 10018, 10018, 10018, 10018, 10046, 10046, 
    10046, 10054, 10054, 10054, 10054, 10121, 10084, 10084, 10084, 10084, 
    10084, 10084, 10084, 10084, 10084, 10084, 10084, 10084, 10084, 10084, 
    10084, 10084, 10084, 10084, 10084, 10084, 9930, 9930, 10084, 10084, 
    10084, 10084, 10084, 10084, 10084, 9930, 9930, 9930, 9930, 9930, 9930,
  9832, 9832, 9580, 8671, 8910, 9103, 8912, 8813, 8981, 8541, 8482, 8514, 
    8469, 8548, 8963, 9449, 9560, 9756, 8887, 9647, 9831, 10015, 10018, 
    10018, 10018, 10018, 10018, 10018, 9849, 9854, 10004, 10018, 10018, 
    10018, 10018, 10018, 10018, 10018, 10018, 10018, 10018, 10018, 10018, 
    10018, 10018, 10012, 10012, 10004, 10014, 10018, 10018, 10046, 10046, 
    10054, 10054, 10054, 10054, 10054, 10054, 10054, 10121, 10084, 10130, 
    10084, 10084, 10084, 10084, 10084, 10084, 10084, 10084, 10084, 10084, 
    10084, 10084, 10084, 10084, 10084, 10084, 10084, 10084, 9930, 9930, 9930, 
    10084, 10084, 10084, 10084, 10084, 9930, 9930, 9930, 9930, 9930, 9930, 
    9930,
  9930, 9832, 9082, 8872, 8653, 9079, 9180, 8906, 9047, 8707, 8567, 8413, 
    8525, 8589, 9249, 9796, 9627, 9714, 9502, 9552, 9939, 10018, 10018, 
    10018, 10018, 10018, 10018, 10018, 10018, 9918, 10018, 10018, 10004, 
    10018, 10018, 10018, 10018, 10018, 10018, 10018, 10018, 10018, 10018, 
    10018, 10018, 9990, 10010, 10018, 10046, 10046, 10046, 10054, 10054, 
    10054, 10054, 10054, 10054, 10054, 10054, 10083, 10084, 10084, 10084, 
    10084, 10084, 10084, 10084, 10084, 10084, 10084, 10084, 10084, 10084, 
    10084, 10084, 10084, 10084, 10084, 10084, 10084, 10084, 9930, 9930, 9930, 
    10084, 10084, 10084, 10084, 10084, 9930, 9930, 9930, 9930, 9930, 9930, 
    9930,
  9880, 9779, 8956, 8945, 8811, 8902, 9182, 9057, 9133, 8786, 8358, 8349, 
    8513, 8294, 9224, 9762, 9529, 9284, 9806, 9831, 9992, 10018, 10018, 
    10018, 10018, 10018, 10018, 10018, 10018, 9990, 9999, 10018, 9976, 10012, 
    10018, 10018, 10018, 9990, 10012, 10012, 10018, 10018, 10018, 10018, 
    9872, 9949, 10043, 10046, 10046, 10054, 10054, 10054, 10054, 10054, 
    10054, 10054, 10054, 10054, 10083, 10083, 10084, 9930, 10084, 10084, 
    10084, 10084, 10084, 10084, 10084, 10084, 10084, 10084, 10084, 10084, 
    10084, 10084, 10084, 10084, 10084, 10084, 10084, 9930, 9930, 10084, 
    10084, 10084, 10084, 10084, 10084, 9930, 9930, 9930, 9930, 9930, 9930, 
    9930,
  9943, 9672, 8863, 8644, 8658, 8979, 9192, 9082, 8998, 8970, 8199, 8627, 
    8725, 8395, 9116, 9629, 9643, 9263, 9668, 9781, 9987, 10018, 10018, 
    10018, 10018, 10018, 10018, 10018, 10018, 10018, 10008, 10018, 10018, 
    9977, 9852, 9864, 9969, 9912, 9836, 9740, 9935, 10018, 10018, 9963, 9884, 
    10008, 10026, 10054, 10054, 10054, 10054, 10054, 10054, 10054, 10054, 
    10054, 10054, 10054, 10107, 10121, 10084, 10084, 10084, 10084, 10084, 
    10084, 10084, 10084, 10084, 10084, 10084, 10084, 10084, 10084, 10084, 
    10084, 10084, 10084, 10084, 10084, 10084, 10084, 10084, 10084, 10084, 
    10084, 10084, 10084, 10084, 9930, 9930, 9930, 9930, 9930, 9930, 9930,
  9990, 9612, 8501, 8432, 8801, 8936, 9230, 9042, 9072, 8954, 8747, 8815, 
    8621, 8638, 8678, 9679, 9619, 9244, 9647, 9974, 9953, 10018, 10018, 
    10018, 10018, 10018, 10018, 10018, 10018, 9976, 10018, 10018, 9976, 9969, 
    9801, 9759, 9864, 9822, 9903, 9598, 9911, 9935, 10046, 10031, 9870, 
    10027, 10054, 10054, 10054, 10054, 10054, 10054, 10054, 10054, 10054, 
    10054, 10054, 10084, 10084, 10084, 10084, 10084, 10084, 10084, 10084, 
    10084, 10084, 10084, 10084, 10084, 10084, 10084, 10084, 10084, 10084, 
    10084, 10084, 10084, 10084, 10084, 10084, 10084, 10084, 10084, 10084, 
    10084, 10084, 10084, 10084, 9930, 9930, 9930, 9930, 9930, 9930, 9930,
  10008, 9544, 8811, 8551, 8877, 9118, 9230, 9067, 9230, 9177, 8815, 8861, 
    8904, 8683, 8979, 9629, 9729, 9680, 9661, 9953, 10018, 10018, 10018, 
    10018, 10018, 10018, 10018, 10018, 10018, 10018, 10025, 10018, 10018, 
    9888, 9966, 9794, 9931, 9918, 9943, 9941, 9992, 10029, 10041, 10054, 
    9915, 10023, 10054, 10054, 10054, 10054, 10083, 10062, 10074, 10054, 
    10054, 10101, 10116, 10084, 10084, 10084, 10084, 10084, 10084, 10084, 
    10084, 10084, 10084, 10084, 10084, 10084, 10084, 10084, 10084, 10084, 
    10084, 10084, 10084, 10084, 10084, 10084, 10084, 10084, 10084, 10084, 
    10084, 10084, 10084, 10084, 9930, 9930, 9930, 9930, 9930, 9930, 9930, 9930,
  9963, 9646, 9019, 8770, 9049, 9021, 8945, 8842, 9005, 9320, 9070, 9173, 
    8919, 8852, 8883, 9634, 9607, 9796, 9706, 9994, 10018, 10018, 10018, 
    10018, 10018, 10018, 10018, 10018, 10018, 9963, 10046, 9963, 10018, 
    10018, 9877, 9894, 9905, 9862, 9930, 9895, 9955, 10046, 10054, 10054, 
    10054, 10054, 10054, 10054, 10083, 10083, 10111, 10102, 10054, 10084, 
    10104, 10084, 10084, 10084, 10084, 10084, 10084, 10084, 10084, 10084, 
    10084, 10084, 10084, 10084, 10084, 10084, 10084, 10084, 10084, 10084, 
    10084, 10084, 10084, 10084, 10084, 10084, 10084, 10084, 10084, 10084, 
    10084, 10084, 10084, 10084, 10084, 9930, 9930, 9930, 9930, 9930, 9930, 
    9930,
  9976, 9296, 8791, 8831, 9067, 9051, 9130, 9065, 9196, 9318, 9422, 9521, 
    8828, 8680, 8770, 9540, 9511, 9695, 9524, 9503, 10002, 10018, 10018, 
    10018, 10012, 10018, 10012, 10018, 10018, 10004, 10007, 10004, 10014, 
    10018, 9920, 9860, 9884, 9842, 9915, 9861, 9925, 10041, 10054, 10054, 
    10054, 10054, 10101, 10083, 10084, 10084, 10121, 10084, 10084, 10084, 
    10084, 10084, 10084, 10084, 10084, 10084, 10084, 10084, 10084, 10084, 
    10084, 10084, 10084, 10084, 10084, 10084, 10084, 10084, 10084, 10084, 
    10084, 10084, 10084, 10084, 10084, 10084, 10084, 10084, 10084, 10084, 
    10084, 10084, 10084, 10084, 10084, 9930, 9930, 9930, 9930, 9930, 9930, 
    9930 ;

 TPW =
  121, 129, 147, 108, 106, 119, 142, 190, 274, 249, 171, 221, 208, 235, 273, 
    285, 309, 255, 200, 184, 219, 255, 247, 273, 269, 286, 272, 247, 256, 
    260, 245, 234, 231, 239, 234, 212, 183, 178, 182, 169, 194, 171, 183, 
    180, 180, 177, 170, 175, 165, 186, 158, 168, 174, 177, 166, 133, 125, 
    121, 118, 99, 111, 116, 110, 101, 94, 91, 96, 91, 94, 95, 100, 93, 90, 
    94, 89, 95, 100, 101, 101, 105, 113, 127, 117, 107, 107, 103, 126, 123, 
    103, 128, 132, 123, 132, 122, 130, 133,
  123, 123, 156, 133, 128, 155, 211, 279, 259, 213, 235, 239, 201, 182, 271, 
    322, 311, 268, 215, 184, 236, 244, 239, 258, 260, 272, 276, 251, 263, 
    256, 227, 206, 206, 194, 202, 196, 180, 188, 186, 190, 210, 184, 186, 
    178, 181, 181, 173, 173, 182, 164, 203, 192, 184, 165, 149, 168, 131, 
    116, 119, 115, 99, 111, 110, 101, 95, 96, 93, 95, 94, 97, 90, 101, 88, 
    94, 89, 93, 100, 106, 109, 123, 121, 122, 115, 106, 102, 102, 96, 118, 
    104, 118, 134, 124, 128, 125, 130, 123,
  157, 161, 173, 158, 192, 269, 283, 288, 197, 260, 183, 205, 177, 248, 264, 
    345, 314, 279, 225, 214, 253, 245, 230, 230, 237, 230, 243, 226, 235, 
    227, 218, 209, 206, 200, 200, 189, 190, 190, 233, 220, 193, 167, 170, 
    187, 186, 189, 190, 183, 178, 153, 192, 181, 183, 175, 147, 150, 137, 
    117, 117, 107, 110, 97, 102, 110, 98, 87, 93, 99, 101, 98, 101, 99, 95, 
    96, 110, 102, 100, 111, 119, 119, 117, 109, 105, 108, 99, 94, 94, 97, 
    118, 107, 127, 123, 133, 127, 130, 130,
  169, 188, 254, 209, 236, 266, 286, 255, 201, 254, 151, 175, 212, 220, 267, 
    299, 295, 298, 246, 256, 252, 262, 242, 237, 245, 251, 241, 241, 212, 
    200, 194, 182, 204, 193, 187, 184, 181, 167, 192, 194, 224, 179, 183, 
    174, 184, 184, 182, 175, 173, 161, 153, 146, 171, 187, 166, 142, 129, 
    128, 122, 105, 108, 92, 99, 101, 93, 92, 96, 102, 103, 101, 95, 90, 104, 
    112, 109, 99, 97, 111, 111, 113, 110, 117, 112, 104, 100, 102, 100, 100, 
    101, 102, 123, 126, 124, 133, 131, 124,
  230, 256, 288, 235, 269, 254, 278, 208, 206, 224, 159, 163, 232, 206, 218, 
    293, 314, 313, 244, 272, 242, 254, 295, 228, 216, 233, 232, 232, 215, 
    225, 193, 212, 198, 188, 195, 190, 191, 191, 182, 176, 188, 195, 178, 
    173, 181, 180, 199, 165, 175, 163, 179, 176, 194, 169, 154, 155, 132, 
    123, 108, 105, 113, 91, 104, 102, 90, 98, 107, 109, 102, 102, 103, 106, 
    123, 123, 116, 111, 105, 110, 107, 109, 108, 84, 82, 89, 103, 109, 100, 
    104, 111, 124, 127, 125, 134, 133, 129, 132,
  302, 332, 314, 273, 230, 268, 279, 188, 237, 174, 213, 273, 243, 220, 263, 
    309, 304, 313, 248, 228, 242, 240, 311, 226, 218, 227, 225, 230, 227, 
    206, 194, 200, 203, 198, 198, 198, 186, 201, 187, 185, 194, 198, 208, 
    184, 185, 217, 212, 183, 165, 192, 195, 196, 147, 135, 128, 126, 115, 
    113, 102, 115, 104, 101, 113, 103, 93, 105, 100, 111, 101, 102, 116, 119, 
    115, 122, 120, 114, 102, 107, 110, 104, 99, 96, 90, 110, 105, 102, 103, 
    100, 94, 126, 125, 120, 130, 125, 132, 136,
  268, 307, 297, 314, 242, 267, 242, 221, 273, 226, 198, 204, 224, 172, 248, 
    310, 293, 216, 235, 253, 279, 243, 220, 207, 211, 208, 208, 204, 206, 
    221, 191, 197, 181, 192, 179, 186, 220, 210, 185, 198, 209, 213, 218, 
    268, 238, 227, 180, 162, 144, 165, 170, 155, 144, 142, 142, 121, 110, 
    107, 110, 108, 103, 88, 101, 98, 111, 108, 95, 102, 101, 113, 118, 122, 
    113, 118, 114, 115, 119, 116, 110, 93, 100, 102, 99, 107, 103, 88, 94, 
    96, 87, 124, 122, 119, 114, 128, 127, 134,
  288, 301, 281, 234, 224, 267, 215, 249, 218, 251, 191, 233, 202, 178, 186, 
    213, 228, 175, 203, 229, 239, 224, 218, 196, 194, 207, 203, 219, 206, 
    200, 194, 202, 206, 185, 185, 184, 207, 197, 203, 210, 222, 297, 283, 
    283, 240, 204, 175, 187, 186, 162, 151, 131, 143, 123, 122, 115, 107, 
    106, 116, 107, 117, 99, 109, 111, 110, 106, 109, 119, 103, 121, 125, 125, 
    111, 126, 123, 117, 126, 117, 113, 106, 98, 96, 99, 102, 97, 99, 99, 101, 
    94, 115, 115, 116, 129, 131, 138, 131,
  259, 375, 201, 171, 203, 191, 213, 319, 259, 229, 211, 215, 170, 180, 146, 
    218, 216, 174, 209, 248, 219, 221, 213, 201, 195, 198, 241, 210, 178, 
    194, 201, 198, 209, 195, 186, 204, 279, 276, 235, 215, 290, 268, 241, 
    212, 191, 181, 139, 153, 137, 134, 129, 156, 136, 118, 134, 109, 111, 
    144, 112, 107, 115, 113, 122, 99, 97, 93, 104, 102, 116, 121, 115, 117, 
    117, 123, 122, 114, 114, 117, 117, 107, 99, 98, 95, 94, 99, 101, 102, 
    111, 100, 120, 121, 118, 122, 127, 131, 138,
  390, 341, 221, 202, 301, 211, 261, 270, 278, 273, 228, 208, 170, 158, 149, 
    201, 200, 216, 188, 205, 199, 213, 197, 212, 196, 196, 199, 192, 200, 
    202, 195, 207, 207, 213, 213, 206, 236, 221, 210, 201, 242, 211, 235, 
    208, 178, 166, 148, 130, 135, 134, 124, 118, 124, 118, 98, 123, 120, 120, 
    118, 114, 111, 117, 113, 106, 108, 108, 96, 113, 121, 119, 122, 123, 114, 
    127, 124, 121, 117, 113, 114, 110, 99, 99, 102, 101, 100, 99, 116, 107, 
    123, 115, 119, 111, 110, 117, 113, 124,
  367, 354, 233, 252, 291, 245, 266, 246, 262, 283, 225, 206, 157, 152, 167, 
    195, 204, 202, 185, 199, 200, 185, 182, 203, 189, 181, 198, 191, 203, 
    204, 208, 206, 197, 221, 207, 228, 220, 206, 215, 199, 218, 213, 226, 
    179, 137, 131, 126, 132, 137, 143, 141, 131, 120, 126, 126, 119, 131, 
    120, 107, 106, 113, 113, 107, 101, 100, 99, 102, 106, 118, 120, 114, 119, 
    121, 124, 116, 114, 105, 109, 122, 106, 95, 97, 106, 94, 98, 109, 101, 
    97, 96, 116, 110, 106, 109, 107, 102, 122,
  345, 300, 220, 248, 244, 292, 218, 214, 287, 250, 226, 212, 183, 142, 147, 
    188, 168, 189, 182, 187, 196, 182, 166, 183, 187, 204, 215, 189, 198, 
    193, 204, 193, 209, 205, 239, 237, 230, 212, 228, 234, 240, 223, 167, 
    142, 137, 135, 133, 126, 103, 99, 123, 108, 103, 105, 116, 111, 117, 117, 
    114, 119, 114, 103, 104, 106, 96, 98, 103, 104, 112, 125, 123, 122, 135, 
    122, 110, 111, 106, 112, 115, 98, 95, 103, 105, 101, 97, 103, 104, 106, 
    106, 122, 111, 100, 99, 96, 103, 118 ;

 TSkin =
  31455, 31334, 30871, 30903, 31094, 31044, 30705, 30574, 29915, 29515, 
    29805, 29656, 29537, 29815, 29982, 29013, 28936, 29112, 29043, 28967, 
    29022, 28762, 28757, 28653, 28683, 28920, 28793, 28852, 28661, 28598, 
    28443, 28256, 27738, 28055, 28031, 27772, 27948, 27450, 27633, 27508, 
    27803, 27856, 27709, 27388, 27649, 27651, 27551, 27674, 27613, 28287, 
    27478, 27691, 27850, 27834, 27766, 27785, 27992, 28078, 27729, 26899, 
    26427, 28260, 28317, 28199, 28160, 28103, 28106, 28104, 28062, 28076, 
    28029, 28048, 28002, 28056, 28108, 28025, 28042, 28067, 28063, 27958, 
    28005, 28057, 27896, 27891, 27941, 27861, 27176, 27343, 27761, 27908, 
    28012, 27657, 27518, 27727, 27822, 27938,
  31374, 31210, 30858, 30733, 30684, 30827, 30330, 29861, 29181, 29797, 
    29437, 29357, 29717, 29690, 29731, 29632, 29386, 29238, 29140, 28956, 
    28855, 28615, 28627, 28343, 28783, 28854, 28837, 28610, 28464, 28539, 
    28543, 28286, 27956, 27993, 27751, 27804, 27786, 27746, 27605, 27922, 
    28004, 27546, 27445, 27644, 27594, 27760, 27861, 27910, 27698, 27646, 
    27739, 27799, 27673, 27841, 27787, 27412, 27191, 27617, 27934, 27210, 
    28271, 28102, 28238, 28208, 28116, 28082, 28068, 27956, 28099, 27974, 
    28004, 27939, 28004, 28073, 28010, 28012, 28099, 28034, 28100, 27990, 
    28039, 28050, 27857, 27933, 27994, 27821, 27765, 27273, 27612, 27595, 
    27572, 27201, 27487, 27656, 27762, 27892,
  31549, 31002, 30729, 30761, 30546, 30276, 30070, 29394, 29871, 29519, 
    29598, 29596, 29685, 29571, 29604, 29828, 29492, 29229, 29085, 29062, 
    28655, 28705, 28754, 28656, 28538, 28459, 28544, 28450, 28622, 28504, 
    28445, 28302, 28240, 27984, 27967, 27845, 27788, 27718, 27488, 27837, 
    27617, 27550, 27693, 27674, 27774, 27845, 27933, 28074, 27831, 27947, 
    27826, 27878, 27901, 27880, 27647, 27549, 27505, 27390, 27410, 27666, 
    27021, 28096, 28033, 28182, 28231, 28133, 28119, 28069, 28024, 27892, 
    27955, 27946, 27990, 28055, 28086, 27958, 28035, 28045, 27988, 27984, 
    27958, 27964, 27920, 27981, 27866, 27670, 27758, 27658, 27172, 27511, 
    27210, 27206, 27583, 27594, 27559, 27792,
  31385, 30818, 30528, 30403, 30253, 30124, 29537, 29449, 29857, 29385, 
    29522, 29614, 29359, 29023, 29449, 29337, 29091, 29492, 29427, 29008, 
    28910, 28505, 28376, 28417, 28491, 28613, 28372, 28332, 28350, 28499, 
    28476, 28281, 28294, 27815, 27672, 27534, 27623, 27511, 27329, 27372, 
    27678, 27696, 27792, 27843, 27924, 28059, 28022, 27992, 28063, 28060, 
    27918, 27920, 27950, 28038, 28005, 27697, 27929, 27811, 27326, 27531, 
    27279, 28083, 28122, 28101, 28136, 28041, 28193, 28075, 27969, 27845, 
    27970, 28056, 28010, 28043, 28060, 27964, 28081, 27905, 27978, 27918, 
    27905, 27560, 27693, 27795, 27895, 27730, 27740, 27593, 27634, 27560, 
    27429, 27356, 27474, 27560, 27567, 27708,
  31032, 30771, 30360, 30348, 30110, 29425, 29199, 29181, 29796, 29554, 
    29624, 29596, 29573, 29082, 29169, 28864, 29624, 29365, 29281, 28749, 
    28730, 27994, 28524, 28232, 28599, 28351, 28232, 28400, 28453, 28682, 
    28342, 28386, 28267, 27909, 28002, 27966, 27884, 27606, 27513, 27585, 
    27803, 27863, 27604, 27932, 28171, 28460, 28197, 28210, 28128, 28139, 
    28175, 28162, 28089, 28081, 28081, 28014, 28041, 27741, 27439, 27731, 
    26963, 28145, 26829, 28207, 28070, 28101, 28093, 27945, 28017, 28069, 
    27944, 28082, 28042, 27903, 28033, 27925, 28079, 28022, 27930, 27888, 
    27826, 26660, 26958, 26991, 27818, 27752, 27664, 27642, 27544, 27215, 
    27451, 27408, 27502, 27564, 27896, 27593,
  30364, 29997, 30339, 30002, 30242, 29614, 28921, 29864, 29767, 29697, 
    29220, 29906, 29397, 29206, 28947, 29279, 29534, 28892, 28788, 28650, 
    28510, 28367, 28633, 28369, 28400, 28382, 28363, 28161, 28456, 28342, 
    28378, 28266, 28218, 28123, 28032, 27933, 27925, 27804, 27841, 27978, 
    27789, 27832, 28005, 28110, 28276, 28476, 28420, 28199, 28020, 28200, 
    28063, 28356, 28255, 28146, 28276, 28266, 28223, 27926, 27773, 27260, 
    28227, 28092, 28033, 28134, 28164, 28145, 28159, 27991, 27908, 27909, 
    27963, 27990, 28008, 28021, 27957, 27973, 28005, 28088, 28077, 27963, 
    27883, 26828, 26771, 26915, 27812, 27658, 27662, 27603, 27494, 27208, 
    27256, 27261, 27280, 27435, 27575, 27638,
  30424, 30649, 30263, 29575, 30006, 29047, 29209, 29889, 29789, 29359, 
    29195, 29351, 29119, 28889, 28891, 29136, 28911, 28869, 28624, 28143, 
    28314, 28340, 28269, 28200, 28303, 28277, 28305, 28121, 28303, 28579, 
    28282, 28236, 27979, 28001, 28009, 28247, 28130, 28110, 28249, 28024, 
    28313, 28162, 28699, 29713, 29235, 28848, 28096, 28292, 27879, 27866, 
    28184, 28457, 28420, 28487, 28108, 28286, 28360, 28188, 27224, 26932, 
    28032, 26508, 28042, 28198, 27915, 27947, 27933, 27902, 27964, 27888, 
    27941, 27902, 27953, 27894, 27904, 27958, 27993, 27867, 27945, 27805, 
    27866, 27050, 27094, 27688, 27678, 27704, 27563, 27544, 27520, 27102, 
    27420, 27352, 27360, 27186, 27524, 27421,
  30204, 30169, 29864, 29764, 28989, 29718, 29983, 29918, 29880, 28740, 
    29123, 29284, 29205, 29089, 28757, 28496, 28711, 28641, 28394, 28539, 
    28443, 27859, 28281, 28329, 28328, 28339, 28095, 28050, 28376, 28462, 
    28270, 28150, 28061, 28102, 28265, 28445, 28291, 28114, 28121, 28436, 
    28661, 29365, 30184, 29993, 28418, 28743, 28534, 28085, 27864, 27917, 
    28069, 28614, 28608, 28486, 28259, 28415, 28302, 27966, 27388, 26926, 
    28000, 28077, 28130, 27960, 28008, 27928, 27825, 27872, 27888, 27911, 
    28023, 27987, 27947, 27884, 27877, 27888, 27877, 27915, 27855, 27936, 
    27880, 27856, 27781, 27680, 27665, 27628, 27628, 27552, 27562, 27385, 
    27275, 27321, 26996, 27161, 27279, 27482,
  30267, 29658, 29847, 29628, 29473, 29995, 29999, 30162, 29489, 29052, 
    29488, 29328, 29337, 28981, 29083, 28690, 28709, 28425, 28464, 28361, 
    27991, 28002, 28282, 28233, 28279, 28256, 27915, 27965, 28247, 28331, 
    28302, 28182, 28035, 28279, 28355, 28395, 29416, 29148, 28536, 28548, 
    29122, 29215, 28421, 28490, 28207, 28153, 27631, 27961, 28072, 28287, 
    28542, 28269, 28475, 28547, 28528, 28104, 27931, 28323, 28150, 28063, 
    28137, 28096, 28022, 28058, 27977, 28020, 27889, 27856, 27952, 28044, 
    28016, 27992, 27879, 27930, 27863, 27969, 27966, 27877, 27835, 27840, 
    27826, 27817, 27767, 27737, 27671, 27773, 27621, 27595, 27569, 27272, 
    27303, 27272, 27028, 27288, 27426, 27492,
  29714, 29773, 29685, 29391, 30359, 29972, 29607, 29024, 29414, 29468, 
    29404, 29231, 28934, 29293, 29156, 28604, 28544, 28504, 28657, 28446, 
    28273, 28315, 28272, 28364, 28359, 28330, 28355, 28236, 28345, 28251, 
    28127, 27983, 28047, 28302, 28304, 28254, 28476, 28025, 28095, 28116, 
    28497, 28400, 28251, 28495, 27860, 27704, 27734, 27950, 27942, 28276, 
    28349, 28391, 28266, 28248, 28177, 27437, 26898, 28093, 28197, 28062, 
    28058, 28063, 28074, 27963, 27959, 27971, 27970, 27979, 27954, 27866, 
    27983, 27830, 27994, 27779, 27902, 27897, 27724, 27764, 27868, 27812, 
    27836, 27717, 27691, 27695, 27691, 27721, 27697, 27547, 27310, 27501, 
    27381, 27182, 27248, 27228, 27204, 27528,
  29646, 29612, 29442, 29689, 30263, 29343, 29188, 29740, 29736, 29559, 
    29506, 29311, 29197, 29073, 29040, 28695, 28666, 28639, 28505, 28347, 
    28334, 28112, 28325, 28452, 28282, 28196, 28427, 28321, 28368, 28165, 
    28045, 28198, 28000, 28360, 28371, 28334, 28612, 28298, 28382, 28529, 
    28483, 28371, 28650, 27760, 27678, 27969, 27901, 27915, 27813, 27758, 
    27549, 27756, 27575, 28264, 26763, 27966, 28115, 28146, 28115, 28091, 
    28110, 28081, 27985, 27933, 27969, 27959, 27925, 28021, 27899, 27936, 
    27874, 27884, 27941, 27797, 27822, 27842, 27881, 27774, 27736, 27729, 
    27729, 27650, 27707, 27697, 27716, 27662, 27722, 27676, 27631, 27493, 
    27347, 27029, 27273, 26875, 27087, 27050,
  29620, 29910, 29223, 29663, 29566, 29081, 30016, 30078, 29740, 29392, 
    29502, 29446, 29161, 29165, 29152, 28726, 28574, 28525, 28529, 28523, 
    28536, 28199, 28430, 28056, 28340, 28369, 28288, 28148, 28033, 28392, 
    28262, 27967, 28093, 28138, 28605, 28658, 28559, 28427, 28280, 28778, 
    28679, 28163, 27876, 27675, 27745, 27853, 27717, 27367, 28440, 28281, 
    27011, 28037, 28100, 28205, 27969, 28055, 28118, 28168, 28174, 28064, 
    27971, 27965, 27923, 27817, 27875, 27868, 27859, 27977, 27910, 27902, 
    27877, 27877, 27837, 27833, 27888, 27883, 27841, 27849, 27793, 27772, 
    27705, 27678, 27718, 27764, 27666, 27682, 27713, 27579, 27563, 27438, 
    27188, 27042, 27092, 26871, 26923, 27031 ;

 WindDir =
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888 ;

 WindSp =
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888 ;

 WindU =
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888 ;

 WindV =
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888 ;

 YM =
  28574, 28517, 27812, 27081, 25757, 24124, 22732, 22208, 22104, 22510, 
    22914, 23625, 24641, 25803, 26662, 28609, 28850, 27869, 27222, 26543, 
    25502, 24375,
  28556, 28508, 27850, 27118, 25897, 24264, 22794, 22228, 22165, 22515, 
    22917, 23480, 24465, 25968, 26713, 28519, 28769, 27769, 27153, 26413, 
    25330, 24241,
  28510, 28484, 27837, 27143, 25951, 24365, 22885, 22307, 22150, 22487, 
    22931, 23394, 24581, 25756, 26676, 28499, 28582, 27588, 26987, 26220, 
    25146, 24134,
  28444, 28449, 27854, 27167, 26031, 24448, 22988, 22331, 22150, 22478, 
    22797, 23570, 24487, 25831, 26897, 28451, 28495, 27495, 26801, 25984, 
    24910, 23967,
  28361, 28397, 27840, 27257, 26151, 24535, 23026, 22372, 22167, 22492, 
    22850, 23588, 24536, 25812, 26685, 28413, 28489, 27372, 26649, 25853, 
    24789, 23947,
  28258, 28309, 27826, 27285, 26196, 24627, 23054, 22395, 22155, 22448, 
    22907, 23580, 24526, 25616, 26725, 28399, 28414, 27170, 26457, 25667, 
    24782, 23919,
  28124, 28165, 27738, 27253, 26234, 24711, 23185, 22407, 22184, 22420, 
    22847, 23438, 24521, 25665, 26637, 28237, 28078, 26823, 26160, 25400, 
    24496, 23892,
  27938, 27958, 27554, 27139, 26210, 24730, 23161, 22495, 22233, 22448, 
    22850, 23453, 24385, 25819, 26334, 28029, 27760, 26347, 25794, 25207, 
    24457, 23778,
  27704, 27701, 27406, 26997, 26147, 24752, 23292, 22506, 22204, 22482, 
    22901, 23422, 24439, 25509, 26503, 27751, 27381, 26174, 25676, 25113, 
    24552, 23939,
  27471, 27443, 27048, 26779, 26044, 24749, 23285, 22553, 22256, 22482, 
    22838, 23526, 24294, 25634, 26462, 27117, 26672, 25864, 25449, 24970, 
    24406, 23831,
  27305, 27251, 26782, 26531, 25951, 24727, 23313, 22600, 22297, 22444, 
    22837, 23455, 24387, 25606, 26806, 26413, 25490, 25308, 25139, 24772, 
    24240, 23871,
  27246, 27177, 26617, 26410, 25910, 24786, 23417, 22617, 22247, 22544, 
    22820, 23571, 24344, 25771, 26765, 25984, 24321, 24818, 24953, 24728, 
    24221, 23724,
  27294, 27221, 26676, 26512, 25967, 24830, 23437, 22587, 22316, 22421, 
    22734, 23370, 24310, 25404, 26503, 26121, 24408, 24897, 25001, 24821, 
    24347, 23737,
  27401, 27330, 26969, 26707, 26035, 24926, 23458, 22699, 22293, 22512, 
    22859, 23383, 24206, 25629, 26513, 26540, 24868, 24976, 25042, 24727, 
    24290, 23863,
  27492, 27423, 27179, 26845, 26198, 24981, 23514, 22734, 22357, 22469, 
    22813, 23415, 24169, 25555, 26410, 26984, 26099, 25539, 25241, 24913, 
    24417, 23863,
  27505, 27437, 27154, 26881, 26235, 24979, 23562, 22740, 22310, 22445, 
    22802, 23405, 24270, 25568, 26522, 27157, 26528, 25848, 25490, 25050, 
    24423, 23949,
  27432, 27359, 27116, 26845, 26257, 25057, 23600, 22787, 22359, 22436, 
    22899, 23347, 24354, 25557, 26507, 27226, 26603, 25869, 25489, 25056, 
    24384, 23809,
  27317, 27232, 27101, 26821, 26247, 25124, 23644, 22789, 22458, 22459, 
    22833, 23265, 24176, 25228, 26454, 27276, 26970, 26064, 25641, 25105, 
    24416, 23762,
  27217, 27119, 26946, 26740, 26226, 25062, 23672, 22816, 22385, 22519, 
    22804, 23399, 24195, 25349, 26267, 27166, 27175, 26301, 25744, 25123, 
    24447, 23895,
  27158, 27061, 26935, 26735, 26195, 25126, 23689, 22842, 22370, 22482, 
    22821, 23432, 24380, 25358, 26522, 27179, 27206, 26367, 25840, 25241, 
    24587, 23854,
  27123, 27052, 27025, 26832, 26244, 25118, 23696, 22836, 22458, 22481, 
    22869, 23340, 24340, 25396, 26490, 27303, 27032, 26287, 25832, 25210, 
    24555, 23941,
  27080, 27061, 27107, 26875, 26260, 25193, 23765, 22912, 22463, 22470, 
    22843, 23277, 24305, 25493, 26723, 27384, 26988, 26244, 25778, 25197, 
    24440, 23887,
  27035, 27068, 27050, 26860, 26304, 25184, 23793, 22909, 22487, 22532, 
    22871, 23393, 24320, 25535, 26526, 27423, 27025, 26294, 25771, 25222, 
    24504, 23847,
  27036, 27072, 27040, 26879, 26289, 25201, 23797, 22926, 22518, 22483, 
    22774, 23301, 24184, 25549, 26642, 27423, 27025, 26229, 25791, 25165, 
    24497, 23853,
  27116, 27099, 27126, 26882, 26303, 25224, 23820, 22974, 22498, 22517, 
    22839, 23395, 24206, 25337, 26701, 27454, 26900, 26243, 25715, 25203, 
    24528, 24014,
  27241, 27171, 27204, 26963, 26392, 25266, 23838, 22982, 22503, 22549, 
    22899, 23309, 24198, 25176, 26554, 27499, 26944, 26235, 25839, 25196, 
    24617, 23919,
  27344, 27275, 27254, 26917, 26379, 25307, 23897, 23038, 22527, 22569, 
    22813, 23415, 24191, 25437, 26596, 27487, 27006, 26257, 25763, 25233, 
    24522, 23899,
  27378, 27353, 27182, 26931, 26366, 25248, 23848, 23032, 22529, 22594, 
    22816, 23286, 24062, 25311, 26501, 27412, 26981, 26243, 25782, 25264, 
    24534, 24059,
  27327, 27340, 27128, 26882, 26332, 25251, 23910, 23020, 22570, 22502, 
    22827, 23341, 24208, 25187, 26206, 27343, 26856, 26164, 25728, 25177, 
    24591, 23992,
  27181, 27210, 27118, 26869, 26288, 25282, 23872, 23094, 22582, 22608, 
    22787, 23349, 24138, 25418, 26435, 27290, 26769, 26126, 25651, 25177, 
    24502, 23992,
  26930, 26972, 26999, 26826, 26288, 25223, 23920, 23075, 22532, 22611, 
    22841, 23282, 24193, 25182, 26451, 27285, 26763, 26156, 25707, 25251, 
    24552, 23965,
  26584, 26643, 26851, 26691, 26263, 25312, 23976, 23066, 22575, 22496, 
    22806, 23331, 24220, 25359, 26613, 27221, 26825, 26243, 25818, 25363, 
    24629, 24058,
  26180, 26236, 26641, 26599, 26185, 25223, 23938, 23122, 22578, 22579, 
    22829, 23318, 24141, 25546, 27059, 27109, 26663, 26154, 25817, 25400, 
    24705, 24038,
  25762, 25790, 26557, 26521, 26114, 25329, 23968, 23099, 22640, 22527, 
    22761, 23259, 24278, 25196, 26399, 26956, 26507, 26069, 25714, 25257, 
    24699, 24138,
  25369, 25384, 26460, 26465, 26119, 25225, 23972, 23131, 22648, 22593, 
    22900, 23249, 24113, 25327, 26551, 26860, 26414, 26018, 25672, 25344, 
    24736, 24098,
  25042, 25093, 26273, 26362, 26051, 25239, 24003, 23131, 22636, 22558, 
    22769, 23322, 24199, 25291, 26525, 26782, 26507, 26141, 25838, 25431, 
    24787, 24285,
  24835, 24944, 26179, 26276, 26048, 25236, 23982, 23116, 22674, 22616, 
    22792, 23381, 24291, 25158, 26287, 26704, 26644, 26235, 25982, 25543, 
    24991, 24245,
  24790, 24906, 26110, 26214, 25956, 25180, 24017, 23142, 22715, 22610, 
    22823, 23386, 24187, 25163, 26164, 26563, 26694, 26314, 25996, 25592, 
    24959, 24345,
  24874, 24924, 26141, 26244, 26010, 25233, 23982, 23163, 22674, 22592, 
    22843, 23309, 24130, 25196, 26322, 26446, 26607, 26256, 26024, 25542, 
    24959, 24499,
  24977, 24937, 26281, 26289, 26032, 25214, 23985, 23192, 22662, 22613, 
    22877, 23398, 24174, 25280, 26578, 26449, 26575, 26350, 26016, 25635, 
    25048, 24458,
  24982, 24885, 26288, 26351, 26076, 25250, 24024, 23172, 22727, 22575, 
    22791, 23380, 24184, 25198, 26646, 26460, 26657, 26278, 25982, 25579, 
    24991, 24432,
  24859, 24746, 26054, 26182, 26090, 25284, 24003, 23210, 22732, 22601, 
    22851, 23286, 24007, 25172, 26362, 26173, 26825, 26328, 25982, 25449, 
    24965, 24365,
  24678, 24564, 25712, 26022, 26016, 25314, 24023, 23186, 22718, 22598, 
    22854, 23413, 24236, 25230, 26324, 25804, 26775, 26256, 25795, 25412, 
    24748, 24311,
  24542, 24428, 25659, 25988, 25956, 25273, 24027, 23172, 22741, 22612, 
    22888, 23403, 23957, 25405, 26484, 25747, 26544, 26162, 25740, 25331, 
    24640, 24117,
  24511, 24393, 25729, 26050, 26013, 25244, 24013, 23207, 22744, 22641, 
    22868, 23314, 24041, 25431, 26279, 25803, 26526, 26046, 25644, 25181, 
    24608, 24157,
  24566, 24440, 25768, 26092, 26035, 25241, 23999, 23216, 22673, 22641, 
    22842, 23278, 24100, 25298, 26460, 25685, 26538, 26075, 25664, 25188, 
    24608, 24084,
  24641, 24511, 25798, 26051, 26010, 25250, 24027, 23177, 22691, 22635, 
    22894, 23319, 24147, 25496, 26332, 25663, 26532, 26089, 25629, 25051, 
    24563, 24123,
  24683, 24568, 25778, 26103, 26021, 25273, 24027, 23183, 22738, 22663, 
    22857, 23446, 24203, 25396, 26615, 25657, 26488, 26017, 25637, 25169, 
    24455, 23937,
  24691, 24608, 25735, 26047, 25979, 25230, 23992, 23201, 22762, 22655, 
    22965, 23342, 24186, 25298, 26901, 25601, 26295, 25916, 25581, 25138, 
    24595, 23996,
  24702, 24645, 25757, 26012, 26001, 25214, 23999, 23192, 22735, 22690, 
    22851, 23377, 24137, 25338, 26615, 25585, 26339, 25837, 25450, 25088, 
    24487, 24030,
  24734, 24688, 25753, 26032, 25984, 25292, 24044, 23210, 22756, 22632, 
    22900, 23309, 24246, 25508, 26535, 25700, 26407, 26060, 25595, 25044, 
    24506, 24050,
  24763, 24715, 25826, 26063, 26045, 25233, 23992, 23210, 22735, 22644, 
    22934, 23301, 24129, 25410, 26188, 25747, 26607, 26249, 25637, 25156, 
    24544, 23950,
  24734, 24687, 25938, 26129, 26047, 25295, 23968, 23207, 22738, 22664, 
    22960, 23428, 24394, 25172, 26532, 25825, 26688, 26204, 25657, 25156, 
    24538, 24070,
  24594, 24568, 25981, 26144, 26042, 25230, 23985, 23237, 22753, 22655, 
    22848, 23385, 24194, 25237, 26634, 25825, 26731, 26328, 25754, 25225, 
    24570, 24171,
  24319, 24344, 25768, 26117, 25941, 25262, 23968, 23189, 22800, 22713, 
    23005, 23299, 24204, 25256, 26465, 25666, 26613, 26435, 25899, 25306, 
    24634, 24077,
  23892, 23978, 25550, 25879, 25939, 25242, 23978, 23198, 22811, 22644, 
    22971, 23405, 24174, 25338, 26537, 25421, 26682, 26610, 26037, 25430, 
    24647, 24064,
  23262, 23387, 25352, 25807, 25878, 25200, 23975, 23184, 22785, 22738, 
    22940, 23352, 24105, 25217, 26445, 25279, 26869, 26710, 26154, 25480, 
    24640, 24137,
  22334, 22477, 25233, 25664, 25867, 25160, 23992, 23181, 22791, 22664, 
    22923, 23373, 24244, 25244, 26641, 25048, 27012, 26754, 26160, 25561, 
    24793, 24084,
  21063, 21237, 24518, 25274, 25681, 25149, 23916, 23160, 22797, 22687, 
    22948, 23376, 24327, 25492, 26409, 24100, 26457, 26668, 26141, 25493, 
    24806, 24104,
  19560, 19799, 23154, 24399, 25300, 25032, 23972, 23190, 22774, 22796, 
    22937, 23368, 24217, 25331, 26615, 22499, 25406, 26596, 26210, 25574, 
    24793, 24178,
  18104, 18414, 22143, 23759, 25040, 24931, 23906, 23193, 22745, 22708, 
    23011, 23421, 24355, 25340, 26448, 21421, 25001, 26567, 26224, 25660, 
    24959, 24238,
  17025, 17373, 21920, 23627, 24954, 24945, 23930, 23181, 22815, 22728, 
    23040, 23373, 24261, 25422, 26967, 21510, 25181, 26632, 26307, 25767, 
    24966, 24312,
  16546, 16889, 22006, 23668, 24980, 24878, 23889, 23214, 22824, 22751, 
    22975, 23323, 24311, 25319, 26494, 21763, 25318, 26589, 26362, 25792, 
    25099, 24345,
  16700, 17011, 21994, 23716, 24969, 24931, 23882, 23146, 22792, 22863, 
    22964, 23366, 24353, 25560, 26574, 21685, 25064, 26582, 26342, 25904, 
    25074, 24412,
  17352, 17615, 22176, 23808, 24995, 24926, 23868, 23196, 22851, 22852, 
    23077, 23510, 24271, 25506, 26540, 21681, 24840, 26509, 26314, 25842, 
    25164, 24373,
  18270, 18476, 22684, 24123, 25089, 24870, 23868, 23161, 22810, 22849, 
    22958, 23434, 24218, 25457, 26489, 22130, 24989, 26553, 26410, 25929, 
    25132, 24480,
  19212, 19371, 23289, 24457, 25195, 24853, 23833, 23135, 22789, 22786, 
    23089, 23417, 24356, 25369, 26494, 22872, 25400, 26597, 26363, 25910, 
    25145, 24527,
  19989, 20136, 23675, 24680, 25287, 24862, 23813, 23161, 22819, 22797, 
    23101, 23455, 24260, 25529, 26540, 23377, 25475, 26589, 26370, 25923, 
    25273, 24514,
  20507, 20681, 23771, 24688, 25307, 24889, 23841, 23135, 22878, 22852, 
    23092, 23440, 24272, 25644, 26654, 23560, 25506, 26590, 26370, 25873, 
    25241, 24594,
  20757, 20979, 23784, 24740, 25264, 24825, 23764, 23138, 22875, 22838, 
    23053, 23438, 24336, 25628, 26729, 23498, 25556, 26582, 26294, 25923, 
    25158, 24487,
  20782, 21048, 23647, 24659, 25250, 24806, 23768, 23118, 22840, 22864, 
    23070, 23499, 24297, 25493, 26723, 23328, 25519, 26575, 26274, 25810, 
    25177, 24668,
  20633, 20925, 23642, 24694, 25202, 24786, 23754, 23144, 22849, 22795, 
    23070, 23484, 24441, 25411, 26514, 23236, 25407, 26496, 26253, 25774, 
    25108, 24528,
  20352, 20647, 23719, 24694, 25219, 24764, 23734, 23089, 22829, 22870, 
    22988, 23477, 24325, 25504, 26479, 23255, 25413, 26496, 26253, 25731, 
    25134, 24568,
  19961, 20243, 23549, 24633, 25182, 24688, 23689, 23086, 22838, 22851, 
    22999, 23416, 24330, 25551, 26725, 23107, 25500, 26467, 26260, 25688, 
    25102, 24522,
  19453, 19726, 23395, 24496, 25159, 24697, 23682, 23077, 22827, 22831, 
    22997, 23546, 24308, 25667, 26321, 22861, 25252, 26395, 26116, 25657, 
    25051, 24589,
  18819, 19091, 23068, 24391, 25082, 24636, 23655, 23072, 22865, 22917, 
    23063, 23536, 24291, 25556, 26729, 22576, 25295, 26403, 26116, 25694, 
    25007, 24435,
  18084, 18342, 22782, 24238, 25042, 24641, 23610, 23031, 22833, 22874, 
    23134, 23475, 24170, 25621, 26544, 22238, 25265, 26424, 26157, 25682, 
    25052, 24663,
  17327, 17549, 22364, 24023, 24942, 24549, 23620, 23066, 22853, 22849, 
    23057, 23430, 24414, 25584, 26575, 21895, 25134, 26432, 26192, 25757, 
    25185, 24637,
  16696, 16878, 22232, 23937, 24942, 24577, 23593, 23058, 22830, 22849, 
    23066, 23552, 24279, 25710, 26631, 21621, 25078, 26454, 26206, 25751, 
    25205, 24677,
  16396, 16559, 22321, 23969, 24939, 24566, 23603, 23022, 22898, 22935, 
    23086, 23407, 24435, 25577, 26721, 21635, 25290, 26454, 26192, 25764, 
    25142, 24550,
  16635, 16795, 22431, 24012, 24962, 24524, 23544, 23032, 22854, 22921, 
    23030, 23590, 24445, 25843, 26646, 21874, 25508, 26396, 26124, 25689, 
    25002, 24417,
  17516, 17660, 22813, 24182, 24957, 24446, 23527, 23076, 22887, 22890, 
    23099, 23555, 24522, 25776, 26774, 22308, 25881, 26339, 26028, 25572, 
    24906, 24404,
  18921, 19019, 23455, 24588, 25063, 24438, 23517, 23032, 22863, 23005, 
    22988, 23540, 24376, 25899, 27010, 23047, 25900, 26310, 25917, 25485, 
    24951, 24311,
  20502, 20537, 24354, 25032, 25160, 24441, 23500, 23015, 22896, 22928, 
    23147, 23545, 24312, 25632, 26784, 23958, 26043, 26260, 25897, 25498, 
    24933, 24271,
  21832, 21823, 24869, 25267, 25203, 24388, 23462, 23033, 22905, 22917, 
    23119, 23586, 24470, 25767, 26829, 24561, 26193, 26246, 25882, 25411, 
    24876, 24404,
  22651, 22632, 24998, 25326, 25201, 24388, 23431, 23039, 22905, 22942, 
    23111, 23627, 24653, 25695, 26823, 24507, 26106, 26253, 25904, 25461, 
    24844, 24338,
  23005, 22996, 25026, 25358, 25195, 24363, 23421, 23025, 22864, 22957, 
    23094, 23630, 24639, 25614, 26668, 24322, 26056, 26260, 25925, 25448, 
    25010, 24352,
  23151, 23145, 25021, 25307, 25149, 24282, 23373, 23025, 22923, 22946, 
    23151, 23541, 24567, 25821, 27057, 24188, 26032, 26196, 25904, 25393, 
    24858, 24299,
  23311, 23294, 25186, 25415, 25164, 24288, 23341, 22969, 22935, 22872, 
    23129, 23724, 24437, 25874, 26734, 24520, 26137, 26182, 25747, 25406, 
    24807, 24272,
  23517, 23495, 25551, 25579, 25153, 24221, 23300, 23010, 22935, 22967, 
    23126, 23689, 24792, 25951, 26528, 25315, 26610, 26196, 25807, 25375, 
    24814, 24226,
  23662, 23666, 25566, 25574, 25087, 24137, 23241, 22925, 22886, 22952, 
    23118, 23730, 24787, 25739, 26826, 25402, 26654, 26182, 25768, 25369, 
    24731, 24113,
  23633, 23683, 25450, 25512, 25010, 24098, 23217, 22961, 22924, 23028, 
    23195, 23704, 24738, 25872, 27212, 24974, 26238, 26175, 25801, 25375, 
    24789, 24193,
  23354, 23405, 25405, 25370, 24939, 24070, 23231, 22946, 22913, 23059, 
    23250, 23804, 24837, 26154, 26993, 24569, 26200, 26103, 25789, 25326, 
    24732, 24133,
  22829, 22775, 25149, 25308, 24859, 23936, 23183, 22968, 22913, 22982, 
    23272, 23832, 24768, 26282, 27023, 23898, 26101, 26118, 25775, 25327, 
    24726, 24234,
  22261, 22043, 25182, 25257, 24816, 23925, 23152, 22891, 22899, 23026, 
    23253, 23733, 24788, 26003, 26863, 23716, 26213, 26118, 25720, 25308, 
    24694, 24114,
  22008, 21710, 25276, 25279, 24673, 23808, 23128, 22906, 22888, 23049, 
    23159, 23923, 24828, 26194, 26941, 23864, 26201, 25909, 25555, 25060, 
    24460, 23948,
  28538, 28503, 27847, 27023, 25764, 24134, 22708, 22189, 22107, 22501, 
    22970, 23665, 24656, 25759, 26631, 28632, 28782, 27810, 27201, 26423, 
    25326, 24259,
  28519, 28492, 27875, 27082, 25869, 24283, 22801, 22244, 22154, 22461, 
    22938, 23695, 24621, 25785, 26501, 28564, 28757, 27729, 27079, 26250, 
    25123, 24226,
  28467, 28466, 27782, 27179, 25995, 24380, 22878, 22259, 22174, 22484, 
    22844, 23634, 24587, 25979, 26699, 28446, 28422, 27464, 26760, 25964, 
    24906, 24005,
  28390, 28423, 27831, 27195, 25998, 24470, 22992, 22327, 22162, 22518, 
    22892, 23670, 24670, 25731, 26728, 28393, 28316, 27247, 26554, 25776, 
    24709, 23725,
  28292, 28353, 27804, 27207, 26038, 24553, 23019, 22382, 22167, 22472, 
    22912, 23540, 24446, 25796, 27021, 28429, 28285, 27103, 26320, 25628, 
    24556, 23918,
  28178, 28235, 27743, 27249, 26129, 24612, 23096, 22420, 22202, 22528, 
    22857, 23525, 24509, 25826, 26534, 28351, 28085, 26750, 26120, 25435, 
    24588, 23931,
  28035, 28057, 27526, 27117, 26106, 24646, 23120, 22473, 22170, 22480, 
    22845, 23451, 24369, 25500, 26638, 28101, 27713, 26410, 25754, 25094, 
    24390, 23677,
  27835, 27818, 27390, 26945, 26072, 24696, 23199, 22479, 22225, 22430, 
    22885, 23496, 24450, 25574, 26504, 27762, 27141, 26000, 25534, 25007, 
    24295, 23744,
  27580, 27532, 27131, 26738, 26032, 24695, 23303, 22543, 22233, 22410, 
    22742, 23488, 24405, 25667, 26606, 27189, 26754, 25863, 25444, 24975, 
    24339, 23696,
  27329, 27250, 26829, 26544, 25882, 24732, 23307, 22543, 22257, 22419, 
    22754, 23374, 24336, 25421, 26632, 26476, 25225, 25098, 25052, 24801, 
    24205, 23683,
  27158, 27052, 26504, 26328, 25810, 24689, 23320, 22589, 22280, 22447, 
    22896, 23399, 24338, 25481, 26182, 25857, 24062, 24630, 24817, 24620, 
    24160, 23616,
  27110, 27006, 26439, 26298, 25837, 24779, 23431, 22633, 22268, 22472, 
    22898, 23462, 24372, 25541, 26654, 25701, 23603, 24528, 24782, 24645, 
    24103, 23675,
  27176, 27107, 26665, 26484, 25937, 24866, 23476, 22642, 22265, 22426, 
    22887, 23391, 24355, 25654, 26576, 26171, 24603, 24953, 25003, 24812, 
    24255, 23755,
  27304, 27271, 27017, 26737, 26065, 24933, 23472, 22665, 22329, 22423, 
    22815, 23408, 24310, 25494, 26712, 26760, 25728, 25472, 25236, 24818, 
    24273, 23748,
  27421, 27398, 27135, 26823, 26182, 24972, 23559, 22718, 22343, 22480, 
    22852, 23418, 24386, 25543, 26557, 27137, 26244, 25631, 25236, 24874, 
    24336, 23821,
  27462, 27429, 27189, 26912, 26268, 25030, 23576, 22735, 22380, 22491, 
    22860, 23398, 24359, 25594, 26731, 27260, 26269, 25638, 25318, 24868, 
    24362, 23814,
  27415, 27369, 27144, 26914, 26248, 25100, 23645, 22765, 22389, 22474, 
    22823, 23471, 24206, 25529, 26554, 27329, 26504, 25709, 25346, 24942, 
    24260, 23880,
  27318, 27259, 27029, 26866, 26248, 25089, 23631, 22808, 22407, 22499, 
    22825, 23478, 24166, 25370, 26529, 27344, 26791, 25918, 25477, 24972, 
    24463, 23827,
  27226, 27149, 27012, 26782, 26245, 25120, 23697, 22841, 22430, 22490, 
    22891, 23395, 24285, 25475, 26554, 27238, 26859, 26120, 25621, 25066, 
    24456, 23867,
  27162, 27069, 26991, 26799, 26207, 25114, 23700, 22873, 22485, 22536, 
    22813, 23389, 24309, 25403, 26560, 27292, 26909, 26264, 25704, 25146, 
    24475, 23933,
  27106, 27023, 27141, 26801, 26251, 25125, 23731, 22899, 22470, 22473, 
    22736, 23321, 24323, 25347, 26617, 27359, 26946, 26285, 25745, 25140, 
    24437, 23899,
  27027, 26991, 27126, 26863, 26296, 25172, 23766, 22940, 22485, 22484, 
    22756, 23379, 24249, 25629, 26935, 27462, 27071, 26401, 25841, 25226, 
    24443, 23825,
  26944, 26964, 27095, 26828, 26307, 25195, 23786, 22949, 22525, 22550, 
    22819, 23358, 24313, 25344, 26663, 27473, 27064, 26385, 25848, 25195, 
    24449, 23825,
  26913, 26955, 27042, 26812, 26276, 25262, 23838, 22937, 22487, 22460, 
    22806, 23335, 24232, 25491, 26595, 27409, 27001, 26307, 25799, 25182, 
    24448, 23851,
  26976, 26990, 27026, 26903, 26353, 25287, 23855, 23019, 22498, 22517, 
    22769, 23342, 24281, 25402, 26553, 27462, 26840, 26170, 25716, 25132, 
    24448, 23871,
  27109, 27083, 27159, 26922, 26360, 25268, 23866, 23028, 22551, 22489, 
    22723, 23314, 24086, 25532, 26509, 27501, 26871, 26191, 25729, 25194, 
    24486, 23865,
  27242, 27205, 27174, 26898, 26356, 25245, 23848, 22989, 22518, 22522, 
    22826, 23378, 24201, 25344, 26560, 27451, 26907, 26169, 25737, 25144, 
    24530, 23844,
  27309, 27286, 27174, 26838, 26316, 25262, 23886, 23028, 22533, 22494, 
    22846, 23314, 24162, 25332, 26478, 27446, 26901, 26249, 25751, 25250, 
    24568, 23871,
  27271, 27260, 27113, 26860, 26307, 25259, 23907, 23042, 22565, 22560, 
    22766, 23326, 24214, 25427, 26616, 27418, 27026, 26256, 25804, 25256, 
    24562, 23884,
  27105, 27106, 27095, 26849, 26373, 25267, 23889, 23057, 22529, 22551, 
    22774, 23298, 24107, 25551, 26388, 27407, 27051, 26328, 25867, 25343, 
    24581, 23997,
  26819, 26850, 26965, 26773, 26307, 25281, 23910, 23054, 22579, 22571, 
    22851, 23283, 24147, 25339, 26618, 27357, 26957, 26363, 25957, 25448, 
    24727, 24043,
  26459, 26524, 26740, 26674, 26229, 25295, 23927, 23095, 22614, 22573, 
    22848, 23313, 24250, 25231, 26479, 27226, 26896, 26392, 25991, 25460, 
    24796, 24063,
  26085, 26149, 26613, 26504, 26189, 25233, 23958, 23112, 22599, 22650, 
    22867, 23455, 24240, 25236, 26424, 27103, 26839, 26356, 26026, 25492, 
    24847, 24116,
  25728, 25756, 26532, 26509, 26151, 25238, 23938, 23103, 22640, 22579, 
    22793, 23409, 24193, 25469, 26279, 27039, 26839, 26443, 26046, 25585, 
    24974, 24390,
  25397, 25405, 26448, 26410, 26109, 25233, 23965, 23115, 22628, 22570, 
    22910, 23371, 24232, 25296, 26606, 26981, 26857, 26443, 26046, 25572, 
    24942, 24336,
  25112, 25154, 26410, 26364, 26101, 25238, 24007, 23165, 22678, 22676, 
    22839, 23379, 24306, 25429, 26320, 26829, 26746, 26378, 26067, 25566, 
    25133, 24437,
  24924, 25021, 26314, 26278, 26049, 25246, 23948, 23162, 22678, 22636, 
    22861, 23307, 24264, 25229, 26441, 26691, 26590, 26225, 25942, 25522, 
    25037, 24376,
  24873, 24979, 26257, 26232, 26014, 25162, 23979, 23165, 22690, 22658, 
    22798, 23287, 24239, 25124, 26629, 26635, 26534, 26182, 25935, 25615, 
    25076, 24403,
  24930, 24981, 26229, 26253, 26003, 25193, 23982, 23153, 22689, 22641, 
    22907, 23294, 24182, 25331, 26551, 26557, 26626, 26290, 25956, 25572, 
    25005, 24450,
  24995, 24972, 26279, 26301, 26082, 25246, 24017, 23168, 22760, 22610, 
    22895, 23403, 24269, 25308, 26620, 26451, 26659, 26247, 25984, 25657, 
    24986, 24456,
  24972, 24904, 26240, 26269, 26091, 25261, 24013, 23214, 22742, 22664, 
    22918, 23330, 24325, 25310, 26454, 26388, 26665, 26218, 25921, 25565, 
    24980, 24516,
  24848, 24773, 25895, 26135, 26010, 25249, 24010, 23220, 22710, 22644, 
    22809, 23355, 24197, 25501, 26729, 26073, 26659, 26269, 25873, 25497, 
    24960, 24362,
  24709, 24641, 25674, 25995, 25976, 25283, 24041, 23214, 22739, 22595, 
    22878, 23286, 24172, 25436, 26579, 25710, 26615, 26225, 25866, 25459, 
    24897, 24389,
  24657, 24587, 25651, 25984, 25969, 25272, 23996, 23202, 22768, 22724, 
    22889, 23266, 24236, 25249, 26543, 25624, 26601, 26247, 25851, 25478, 
    24941, 24456,
  24725, 24639, 25737, 26067, 26014, 25269, 24027, 23214, 22727, 22666, 
    22915, 23416, 24162, 25277, 26225, 25685, 26590, 26182, 25804, 25416, 
    24820, 24349,
  24856, 24748, 25920, 26126, 26069, 25291, 24003, 23235, 22745, 22623, 
    22809, 23317, 24271, 25184, 26132, 25835, 26646, 26189, 25790, 25322, 
    24833, 24249,
  24953, 24841, 26160, 26229, 26095, 25280, 24034, 23197, 22794, 22626, 
    22935, 23322, 24224, 25140, 26045, 25925, 26682, 26160, 25728, 25297, 
    24648, 24208,
  24958, 24878, 26085, 26210, 26095, 25238, 24044, 23205, 22788, 22732, 
    22866, 23380, 24115, 25366, 26598, 25928, 26782, 26182, 25735, 25210, 
    24712, 24095,
  24895, 24865, 25793, 26035, 26046, 25286, 24037, 23202, 22745, 22660, 
    22929, 23347, 24204, 25217, 26532, 25704, 26621, 26168, 25707, 25254, 
    24655, 24108,
  24836, 24832, 25719, 26035, 25991, 25243, 24024, 23238, 22741, 22704, 
    22832, 23357, 24061, 25305, 26268, 25549, 26565, 26269, 25700, 25136, 
    24610, 24055,
  24834, 24809, 25726, 26082, 26029, 25277, 24041, 23223, 22771, 22741, 
    22887, 23380, 24157, 25263, 26506, 25591, 26682, 26297, 25721, 25130, 
    24527, 24102,
  24865, 24797, 25801, 26075, 26066, 25283, 24037, 23232, 22841, 22709, 
    22978, 23481, 24194, 25343, 26494, 25624, 26682, 26348, 25756, 25260, 
    24566, 24068,
  24846, 24757, 25849, 26116, 26046, 25254, 24058, 23241, 22815, 22675, 
    22958, 23340, 24182, 25368, 26623, 25682, 26707, 26369, 25845, 25341, 
    24604, 24068,
  24701, 24645, 25857, 26137, 26020, 25283, 23996, 23200, 22797, 22655, 
    22847, 23421, 24236, 25326, 26244, 25769, 26665, 26326, 25851, 25322, 
    24680, 24289,
  24413, 24434, 25788, 26070, 26017, 25229, 23989, 23226, 22809, 22684, 
    22998, 23406, 24337, 25219, 26775, 25644, 26540, 26319, 25804, 25310, 
    24642, 24095,
  24003, 24101, 25387, 25806, 25900, 25196, 24017, 23244, 22771, 22741, 
    22924, 23391, 24251, 25375, 26751, 25270, 26496, 26348, 25859, 25316, 
    24630, 24135,
  23450, 23586, 24926, 25499, 25717, 25216, 23972, 23197, 22780, 22721, 
    22938, 23447, 24207, 25289, 26378, 24786, 26179, 26442, 25970, 25391, 
    24706, 24149,
  22658, 22802, 24924, 25510, 25791, 25137, 23992, 23191, 22856, 22779, 
    22978, 23317, 24251, 25156, 26657, 24749, 26347, 26594, 26073, 25497, 
    24763, 24162,
  21535, 21711, 25007, 25561, 25766, 25126, 23958, 23200, 22842, 22667, 
    22970, 23459, 24261, 25324, 26385, 24813, 26807, 26666, 26107, 25503, 
    24833, 24323,
  20138, 20396, 24188, 25090, 25554, 25109, 23944, 23236, 22833, 22748, 
    22998, 23368, 24301, 25352, 26222, 23727, 26216, 26659, 26212, 25701, 
    24834, 24223,
  18718, 19074, 22916, 24237, 25239, 25003, 23909, 23174, 22807, 22765, 
    23024, 23419, 24247, 25345, 26460, 22228, 25202, 26551, 26335, 25782, 
    24974, 24357,
  17624, 18044, 22079, 23742, 24990, 24911, 23903, 23197, 22780, 22851, 
    22967, 23363, 24210, 25399, 26470, 21527, 25028, 26529, 26315, 25826, 
    25025, 24437,
  17127, 17561, 22046, 23724, 24950, 24860, 23878, 23212, 22842, 22808, 
    23039, 23505, 24144, 25548, 26359, 21754, 25190, 26565, 26309, 25807, 
    25076, 24390,
  17296, 17701, 22412, 23906, 24996, 24911, 23844, 23180, 22837, 22808, 
    22982, 23412, 24321, 25620, 26468, 21930, 25215, 26551, 26350, 25871, 
    25165, 24484,
  17986, 18326, 22625, 24060, 25039, 24902, 23847, 23174, 22810, 22782, 
    23010, 23414, 24265, 25476, 26623, 22130, 25078, 26507, 26295, 25851, 
    25114, 24477,
  18924, 19174, 23102, 24391, 25176, 24911, 23869, 23151, 22843, 22834, 
    23090, 23521, 24205, 25453, 26749, 22675, 25308, 26529, 26343, 25876, 
    25217, 24537,
  19825, 20002, 23649, 24620, 25242, 24852, 23816, 23160, 22817, 22837, 
    23016, 23427, 24240, 25539, 26616, 23321, 25514, 26623, 26357, 25896, 
    25160, 24544,
  20508, 20668, 23862, 24803, 25277, 24866, 23865, 23148, 22813, 22789, 
    23090, 23417, 24285, 25509, 27038, 23649, 25558, 26579, 26344, 25926, 
    25236, 24685,
  20932, 21118, 23931, 24765, 25325, 24872, 23778, 23157, 22864, 22887, 
    23054, 23499, 24463, 25486, 26429, 23635, 25589, 26573, 26316, 26001, 
    25275, 24658,
  21144, 21354, 23746, 24693, 25237, 24821, 23807, 23131, 22843, 22809, 
    23017, 23451, 24251, 25355, 26534, 23518, 25421, 26529, 26310, 25909, 
    25224, 24719,
  21206, 21415, 23792, 24696, 25308, 24796, 23719, 23131, 22861, 22875, 
    23080, 23504, 24217, 25376, 26563, 23459, 25371, 26451, 26241, 25810, 
    25141, 24585,
  21148, 21352, 23936, 24814, 25243, 24797, 23734, 23190, 22847, 22867, 
    23120, 23507, 24236, 25591, 26731, 23567, 25571, 26465, 26192, 25760, 
    25053, 24566,
  20976, 21192, 24018, 24822, 25292, 24721, 23738, 23102, 22859, 22864, 
    23058, 23513, 24337, 25610, 26895, 23670, 25508, 26466, 26157, 25692, 
    25097, 24439,
  20675, 20923, 23919, 24791, 25243, 24727, 23717, 23185, 22867, 22856, 
    23012, 23495, 24370, 25675, 26604, 23575, 25639, 26479, 26172, 25779, 
    25136, 24573,
  20217, 20499, 23792, 24739, 25206, 24710, 23696, 23120, 22874, 22848, 
    23152, 23467, 24523, 25666, 26689, 23413, 25472, 26365, 26103, 25749, 
    25110, 24613,
  19584, 19876, 23516, 24584, 25140, 24699, 23696, 23132, 22853, 22879, 
    23050, 23536, 24338, 25607, 26765, 23156, 25466, 26445, 26157, 25749, 
    25213, 24687,
  18794, 19062, 23119, 24393, 25089, 24696, 23676, 23032, 22880, 22882, 
    23124, 23597, 24425, 25463, 26260, 22763, 25466, 26451, 26151, 25810, 
    25168, 24594,
  17923, 18154, 22713, 24207, 24989, 24539, 23620, 23062, 22868, 22880, 
    23033, 23531, 24423, 25838, 26937, 22313, 25416, 26423, 26159, 25835, 
    25277, 24721,
  17141, 17349, 22427, 24017, 24995, 24562, 23568, 23062, 22904, 22909, 
    23073, 23579, 24400, 25660, 26754, 21981, 25373, 26429, 26151, 25810, 
    25258, 24701,
  16696, 16901, 22359, 24001, 24952, 24554, 23579, 23057, 22851, 22924, 
    23119, 23529, 24512, 25801, 27004, 21914, 25646, 26429, 26132, 25718, 
    25169, 24648,
  16842, 17035, 22486, 24100, 24966, 24493, 23520, 23028, 22820, 22921, 
    23122, 23669, 24460, 25645, 26671, 22066, 25671, 26351, 25979, 25626, 
    24966, 24474,
  17684, 17834, 22798, 24264, 24952, 24484, 23531, 23063, 22884, 22869, 
    23082, 23636, 24312, 25643, 26704, 22361, 25765, 26323, 25946, 25570, 
    24966, 24448,
  19075, 19163, 23563, 24606, 25033, 24420, 23528, 23019, 22870, 22899, 
    23151, 23513, 24495, 25690, 27149, 23105, 25857, 26244, 25932, 25464, 
    24954, 24388,
  20636, 20674, 24399, 25083, 25113, 24406, 23465, 23025, 22905, 22939, 
    23077, 23581, 24375, 25648, 26629, 24045, 26064, 26244, 25857, 25452, 
    24871, 24402,
  21940, 21954, 24947, 25306, 25191, 24370, 23431, 23029, 22897, 22919, 
    23126, 23690, 24649, 25674, 26795, 24627, 26195, 26273, 25906, 25502, 
    24923, 24536,
  22739, 22743, 25071, 25384, 25159, 24351, 23400, 23002, 22897, 22925, 
    23115, 23640, 24671, 25776, 26857, 24596, 26114, 26229, 25926, 25533, 
    25043, 24369,
  23075, 23066, 25066, 25344, 25162, 24317, 23365, 23011, 22865, 22945, 
    23118, 23752, 24605, 25872, 26984, 24490, 26046, 26310, 25960, 25533, 
    24987, 24516,
  23188, 23160, 25087, 25341, 25102, 24292, 23373, 23020, 22915, 22983, 
    23204, 23633, 24464, 25821, 27049, 24364, 26034, 26223, 25844, 25453, 
    24898, 24450,
  23295, 23256, 25067, 25355, 25091, 24245, 23311, 22944, 22889, 22972, 
    23122, 23813, 24689, 25904, 26932, 24464, 26065, 26179, 25831, 25541, 
    24924, 24377,
  23458, 23428, 25244, 25417, 25088, 24186, 23300, 22938, 22877, 22972, 
    23187, 23600, 24729, 25863, 26934, 24879, 26257, 26085, 25700, 25355, 
    24708, 24270,
  23616, 23622, 25341, 25449, 25017, 24156, 23210, 22947, 22936, 22958, 
    23125, 23657, 24682, 25989, 27074, 24882, 26239, 26057, 25769, 25342, 
    24778, 24351,
  23678, 23724, 25265, 25390, 24968, 24069, 23217, 22966, 22863, 22952, 
    23182, 23745, 24567, 25889, 27142, 24594, 26015, 26044, 25694, 25343, 
    24765, 24204,
  23539, 23574, 25298, 25396, 24923, 24008, 23235, 22960, 22913, 22985, 
    23231, 23707, 24697, 26122, 26921, 24479, 26097, 26015, 25694, 25237, 
    24759, 24218,
  23148, 23077, 25315, 25358, 24806, 23960, 23141, 22931, 22911, 22996, 
    23174, 23829, 24813, 26101, 26844, 24158, 26103, 26059, 25653, 25306, 
    24639, 24132,
  22665, 22444, 25263, 25351, 24817, 23885, 23131, 22948, 22897, 22925, 
    23257, 23913, 24880, 26048, 27204, 24054, 26184, 26051, 25715, 25312, 
    24697, 24232,
  22440, 22146, 25346, 25281, 24752, 23809, 23062, 22905, 22943, 23051, 
    23277, 23863, 24794, 26069, 27169, 24039, 26116, 26007, 25584, 25170, 
    24583, 23946,
  28481, 28432, 27793, 27082, 25788, 24139, 22730, 22179, 22165, 22489, 
    22912, 23714, 24769, 25890, 26542, 28678, 28703, 27544, 26949, 26245, 
    25127, 24066,
  28459, 28422, 27804, 27119, 25831, 24276, 22795, 22232, 22127, 22512, 
    22929, 23503, 24559, 25751, 26757, 28535, 28534, 27407, 26701, 25960, 
    24898, 23899,
  28398, 28395, 27699, 27073, 25929, 24371, 22906, 22265, 22173, 22457, 
    22914, 23620, 24643, 25626, 26573, 28443, 28229, 27110, 26363, 25642, 
    24625, 23746,
  28311, 28352, 27747, 27121, 26056, 24461, 22969, 22353, 22178, 22517, 
    22942, 23518, 24539, 25757, 26765, 28310, 28062, 26923, 26156, 25450, 
    24504, 23679,
  28207, 28268, 27656, 27121, 26042, 24519, 23013, 22349, 22178, 22499, 
    22925, 23394, 24487, 25747, 26535, 28306, 27863, 26642, 25888, 25356, 
    24465, 23845,
  28091, 28121, 27582, 27095, 25999, 24581, 23082, 22370, 22137, 22433, 
    22851, 23599, 24440, 25698, 26563, 28132, 27539, 26246, 25673, 25095, 
    24421, 23764,
  27944, 27910, 27415, 26989, 26060, 24614, 23138, 22452, 22245, 22504, 
    22822, 23459, 24425, 25759, 26842, 27848, 27234, 26051, 25508, 24977, 
    24331, 23738,
  27735, 27651, 27194, 26787, 25964, 24637, 23190, 22490, 22218, 22490, 
    22859, 23507, 24361, 25910, 26760, 27368, 26687, 25863, 25467, 24983, 
    24357, 23777,
  27468, 27361, 26842, 26535, 25850, 24667, 23262, 22501, 22268, 22573, 
    22861, 23435, 24513, 25807, 26696, 26607, 25978, 25603, 25315, 24915, 
    24293, 23757,
  27209, 27083, 26447, 26265, 25772, 24681, 23293, 22545, 22268, 22463, 
    22898, 23473, 24385, 25604, 26703, 25924, 24057, 24594, 24784, 24653, 
    24235, 23816,
  27041, 26897, 26403, 26176, 25751, 24717, 23377, 22589, 22311, 22457, 
    22890, 23496, 24485, 25495, 26774, 25659, 24287, 24896, 24963, 24696, 
    24216, 23730,
  27007, 26874, 26501, 26276, 25818, 24784, 23411, 22610, 22308, 22483, 
    22898, 23526, 24391, 25567, 26490, 25941, 24311, 24810, 24893, 24640, 
    24196, 23723,
  27086, 27008, 26657, 26540, 25978, 24876, 23445, 22680, 22302, 22477, 
    22997, 23376, 24386, 25472, 26698, 26472, 25349, 25271, 25128, 24789, 
    24285, 23922,
  27225, 27202, 26981, 26723, 26051, 24899, 23487, 22706, 22340, 22519, 
    22840, 23353, 24388, 25562, 26245, 26975, 26251, 25689, 25293, 24863, 
    24310, 23802,
  27355, 27350, 27059, 26776, 26104, 24949, 23497, 22750, 22354, 22499, 
    22871, 23383, 24309, 25355, 26594, 27176, 26294, 25552, 25203, 24751, 
    24252, 23835,
  27419, 27400, 27125, 26838, 26192, 24988, 23559, 22779, 22386, 22496, 
    22902, 23386, 24178, 25481, 26594, 27304, 26064, 25501, 25175, 24831, 
    24246, 23768,
  27397, 27366, 27157, 26826, 26263, 25010, 23597, 22791, 22424, 22482, 
    22870, 23418, 24361, 25625, 26528, 27346, 26431, 25696, 25327, 24893, 
    24442, 23860,
  27315, 27283, 27076, 26829, 26166, 25120, 23601, 22814, 22452, 22559, 
    22850, 23451, 24193, 25403, 26744, 27351, 26660, 25882, 25471, 24980, 
    24360, 23834,
  27219, 27179, 26991, 26785, 26226, 25100, 23653, 22885, 22438, 22521, 
    22770, 23382, 24180, 25589, 26567, 27310, 26704, 26084, 25560, 25036, 
    24442, 23907,
  27132, 27073, 27075, 26835, 26203, 25122, 23725, 22896, 22463, 22635, 
    22833, 23385, 24380, 25519, 26726, 27301, 26916, 26149, 25663, 25129, 
    24435, 23880,
  27040, 26971, 27072, 26824, 26243, 25158, 23760, 22920, 22437, 22549, 
    22904, 23384, 24335, 25538, 26685, 27378, 27009, 26344, 25850, 25222, 
    24562, 23913,
  26927, 26878, 27026, 26795, 26246, 25110, 23752, 22919, 22504, 22534, 
    22909, 23387, 24246, 25563, 26753, 27400, 27009, 26379, 25870, 25396, 
    24536, 23873,
  26813, 26805, 26957, 26800, 26263, 25136, 23780, 22913, 22545, 22577, 
    22801, 23336, 24216, 25468, 26426, 27378, 27015, 26351, 25815, 25271, 
    24498, 23939,
  26758, 26779, 26922, 26807, 26271, 25217, 23797, 22957, 22515, 22626, 
    22886, 23371, 24117, 25663, 26416, 27406, 27065, 26373, 25849, 25265, 
    24523, 23865,
  26807, 26825, 27041, 26837, 26279, 25208, 23835, 22981, 22553, 22591, 
    22945, 23381, 24389, 25410, 26554, 27439, 27132, 26407, 25959, 25283, 
    24580, 23918,
  26945, 26941, 27099, 26921, 26301, 25233, 23856, 23001, 22542, 22557, 
    22882, 23363, 24164, 25314, 26472, 27498, 27096, 26451, 25945, 25295, 
    24554, 24005,
  27104, 27082, 27148, 26829, 26328, 25214, 23897, 23021, 22559, 22599, 
    22888, 23396, 24205, 25376, 26668, 27398, 26990, 26407, 25951, 25376, 
    24668, 23938,
  27204, 27172, 27107, 26837, 26265, 25247, 23877, 22992, 22561, 22573, 
    22871, 23380, 24188, 25425, 26360, 27389, 26996, 26451, 25979, 25444, 
    24713, 23971,
  27187, 27143, 27104, 26896, 26354, 25292, 23870, 23051, 22605, 22576, 
    22879, 23319, 24232, 25437, 26306, 27437, 27170, 26487, 26013, 25494, 
    24700, 24071,
  27026, 26981, 27010, 26872, 26307, 25272, 23963, 23039, 22634, 22556, 
    22813, 23337, 24126, 25353, 26354, 27409, 27207, 26523, 26076, 25456, 
    24776, 24137,
  26742, 26721, 26950, 26779, 26288, 25261, 23946, 23095, 22625, 22558, 
    22802, 23344, 24128, 25271, 26597, 27365, 27195, 26537, 26082, 25562, 
    24890, 24285,
  26405, 26415, 26747, 26701, 26228, 25294, 23973, 23065, 22651, 22572, 
    22913, 23425, 24215, 25404, 26767, 27275, 27151, 26609, 26172, 25704, 
    24966, 24337,
  26076, 26089, 26635, 26551, 26176, 25289, 23945, 23124, 22640, 22575, 
    22841, 23306, 24303, 25148, 26437, 27129, 27032, 26507, 26157, 25685, 
    24922, 24358,
  25769, 25757, 26556, 26538, 26191, 25238, 23983, 23138, 22657, 22610, 
    22893, 23382, 24133, 25292, 26366, 27066, 26884, 26501, 26137, 25810, 
    25144, 24498,
  25473, 25451, 26470, 26504, 26139, 25221, 23976, 23129, 22674, 22583, 
    22861, 23277, 24172, 25236, 26291, 26979, 26896, 26450, 26165, 25648, 
    25132, 24518,
  25202, 25211, 26384, 26419, 26087, 25241, 24004, 23177, 22706, 22672, 
    22855, 23305, 24137, 25445, 26391, 26841, 26914, 26479, 26151, 25773, 
    25144, 24631,
  25012, 25059, 26237, 26312, 26042, 25215, 23973, 23158, 22703, 22635, 
    22878, 23338, 24212, 25262, 26459, 26666, 26678, 26298, 26075, 25679, 
    25157, 24550,
  24945, 24986, 26201, 26225, 26010, 25179, 23959, 23168, 22671, 22583, 
    22803, 23290, 24204, 25259, 26391, 26554, 26541, 26219, 25874, 25567, 
    25106, 24584,
  24975, 24961, 26135, 26188, 25984, 25196, 24004, 23188, 22697, 22597, 
    22883, 23450, 24053, 25070, 26138, 26429, 26491, 26096, 25819, 25492, 
    25016, 24517,
  25012, 24941, 26188, 26234, 26001, 25215, 23917, 23120, 22732, 22620, 
    22886, 23330, 24081, 25206, 26382, 26390, 26460, 26118, 25771, 25455, 
    25074, 24537,
  24974, 24886, 26049, 26131, 26039, 25226, 23996, 23173, 22715, 22594, 
    22852, 23259, 24179, 25310, 26862, 26192, 26559, 26219, 25840, 25511, 
    25067, 24624,
  24867, 24800, 25823, 26107, 25941, 25221, 23979, 23132, 22762, 22640, 
    22917, 23333, 24258, 25264, 26665, 25872, 26404, 26132, 25819, 25436, 
    24997, 24476,
  24786, 24748, 25782, 26069, 26024, 25246, 24000, 23155, 22732, 22660, 
    22860, 23307, 24181, 25359, 26043, 25763, 26454, 26125, 25819, 25442, 
    24895, 24517,
  24830, 24802, 25949, 26147, 26021, 25229, 24031, 23226, 22738, 22588, 
    22803, 23292, 24073, 25312, 26590, 25832, 26653, 26204, 25832, 25454, 
    24952, 24416,
  25004, 24962, 25954, 26212, 26021, 25285, 23993, 23182, 22714, 22648, 
    22852, 23376, 24097, 25264, 26269, 25876, 26707, 26262, 25901, 25417, 
    24959, 24510,
  25215, 25149, 26074, 26266, 26078, 25282, 24038, 23202, 22773, 22665, 
    22866, 23370, 24132, 25163, 26751, 25928, 26728, 26218, 25819, 25411, 
    24895, 24483,
  25344, 25278, 26301, 26344, 26124, 25268, 24007, 23238, 22750, 22694, 
    22934, 23325, 24219, 25334, 26382, 26179, 26776, 26232, 25776, 25361, 
    24825, 24403,
  25334, 25312, 26272, 26284, 26157, 25263, 24035, 23205, 22782, 22714, 
    22792, 23320, 24055, 25163, 26454, 26192, 26782, 26218, 25764, 25336, 
    24768, 24342,
  25230, 25268, 26157, 26247, 26087, 25254, 24024, 23235, 22767, 22677, 
    22940, 23370, 24272, 25100, 26307, 26003, 26734, 26232, 25750, 25268, 
    24742, 24202,
  25133, 25193, 26031, 26176, 26092, 25243, 23982, 23223, 22773, 22703, 
    22945, 23292, 24184, 25503, 26679, 25854, 26678, 26298, 25729, 25131, 
    24608, 24162,
  25111, 25131, 26010, 26163, 26015, 25263, 23975, 23231, 22805, 22668, 
    22923, 23381, 24191, 25247, 26747, 25875, 26715, 26282, 25701, 25230, 
    24685, 24142,
  25139, 25094, 25960, 26157, 26087, 25251, 24011, 23247, 22832, 22706, 
    22929, 23381, 24327, 25447, 26354, 25829, 26757, 26399, 25867, 25224, 
    24615, 24109,
  25117, 25048, 26064, 26228, 26078, 25296, 24017, 23235, 22838, 22706, 
    22948, 23360, 24300, 25483, 26796, 25847, 26740, 26414, 25888, 25255, 
    24679, 24243,
  24958, 24930, 26020, 26228, 26056, 25207, 23979, 23202, 22794, 22680, 
    22872, 23424, 24083, 25368, 26610, 25900, 26690, 26385, 25840, 25268, 
    24685, 24002,
  24649, 24702, 25857, 26118, 25995, 25232, 24024, 23185, 22797, 22678, 
    22920, 23370, 24196, 25229, 26257, 25726, 26422, 26197, 25688, 25206, 
    24558, 24176,
  24236, 24353, 25506, 25897, 25907, 25212, 23962, 23250, 22756, 22720, 
    22958, 23325, 24298, 25298, 26262, 25320, 26447, 26326, 25819, 25318, 
    24602, 24096,
  23722, 23855, 25070, 25638, 25795, 25117, 23931, 23182, 22788, 22692, 
    22972, 23467, 24103, 25280, 26557, 24766, 26366, 26464, 25971, 25392, 
    24666, 24122,
  23021, 23148, 24958, 25530, 25769, 25128, 23941, 23208, 22794, 22740, 
    22961, 23277, 24196, 25338, 26665, 24643, 26142, 26507, 26081, 25492, 
    24743, 24116,
  22021, 22181, 25047, 25555, 25735, 25181, 24011, 23206, 22821, 22747, 
    22898, 23396, 24143, 25375, 26707, 24894, 26559, 26681, 26206, 25579, 
    24813, 24250,
  20743, 20994, 24720, 25366, 25701, 25117, 23969, 23229, 22847, 22792, 
    22975, 23445, 24103, 25266, 26393, 24529, 26535, 26760, 26248, 25654, 
    24921, 24424,
  19410, 19770, 23617, 24640, 25366, 25061, 23945, 23188, 22827, 22787, 
    23009, 23287, 24389, 25269, 26223, 23206, 25900, 26645, 26275, 25748, 
    25004, 24337,
  18367, 18801, 22535, 23940, 25120, 24952, 23914, 23221, 22844, 22793, 
    22915, 23361, 24306, 25369, 26269, 21967, 24947, 26363, 26268, 25760, 
    24966, 24263,
  17902, 18355, 22383, 23808, 25011, 24887, 23872, 23232, 22821, 22764, 
    23030, 23389, 24256, 25329, 26535, 21950, 25054, 26435, 26289, 25804, 
    25036, 24270,
  18092, 18514, 22725, 24120, 25097, 24896, 23886, 23180, 22833, 22796, 
    22930, 23471, 24247, 25474, 26668, 22401, 25458, 26501, 26275, 25841, 
    25049, 24324,
  18781, 19126, 23037, 24288, 25166, 24843, 23844, 23171, 22827, 22736, 
    22953, 23334, 24133, 25406, 25959, 22701, 25402, 26523, 26303, 25854, 
    25081, 24418,
  19668, 19911, 23503, 24597, 25220, 24899, 23858, 23150, 22836, 22753, 
    22922, 23446, 24148, 25271, 26425, 23093, 25321, 26559, 26338, 25941, 
    25183, 24485,
  20467, 20634, 24001, 24896, 25358, 24919, 23817, 23177, 22816, 22774, 
    22942, 23359, 24279, 25153, 26682, 23722, 25670, 26545, 26351, 25935, 
    25209, 24552,
  21026, 21185, 24132, 24913, 25352, 24846, 23797, 23133, 22836, 22817, 
    22950, 23344, 24247, 25460, 26426, 23911, 25776, 26538, 26359, 25842, 
    25247, 24505,
  21350, 21540, 24051, 24896, 25298, 24855, 23807, 23175, 22880, 22791, 
    22979, 23340, 24299, 25241, 26748, 23800, 25657, 26531, 26276, 25873, 
    25203, 24646,
  21522, 21716, 23978, 24824, 25281, 24815, 23772, 23145, 22790, 22840, 
    22968, 23381, 24245, 25449, 26612, 23657, 25533, 26509, 26269, 25724, 
    25139, 24566,
  21599, 21757, 24088, 24878, 25295, 24841, 23728, 23140, 22869, 22860, 
    23019, 23401, 24302, 25388, 26797, 23754, 25601, 26466, 26187, 25712, 
    25038, 24453,
  21592, 21718, 24275, 24972, 25312, 24768, 23779, 23149, 22849, 22821, 
    22988, 23475, 24231, 25582, 26610, 23885, 25664, 26437, 26179, 25724, 
    25089, 24567,
  21485, 21627, 24235, 24940, 25330, 24732, 23745, 23087, 22840, 22789, 
    23071, 23482, 24298, 25533, 26729, 23935, 25632, 26415, 26179, 25656, 
    24994, 24573,
  21251, 21449, 24154, 24956, 25290, 24760, 23714, 23087, 22885, 22864, 
    23014, 23475, 24434, 25444, 26604, 23912, 25701, 26437, 26132, 25719, 
    25045, 24553,
  20854, 21108, 23997, 24800, 25224, 24701, 23666, 23067, 22885, 22838, 
    23041, 23508, 24367, 25451, 26739, 23800, 25889, 26437, 26076, 25694, 
    25096, 24600,
  20265, 20539, 23863, 24728, 25159, 24659, 23638, 23073, 22847, 22836, 
    23069, 23443, 24406, 25594, 27110, 23632, 25776, 26459, 26146, 25825, 
    25249, 24681,
  19485, 19742, 23480, 24534, 25093, 24626, 23614, 23076, 22870, 22865, 
    23049, 23491, 24370, 25666, 26782, 23211, 25616, 26467, 26132, 25676, 
    25109, 24621,
  18579, 18811, 22999, 24262, 25021, 24556, 23607, 23085, 22853, 22908, 
    23027, 23499, 24392, 25550, 26472, 22690, 25616, 26467, 26167, 25769, 
    25199, 24702,
  17716, 17942, 22543, 24072, 24939, 24542, 23590, 23068, 22898, 22914, 
    23113, 23547, 24366, 25573, 26899, 22235, 25554, 26381, 26112, 25732, 
    25135, 24629,
  17172, 17396, 22414, 24013, 24967, 24565, 23584, 23083, 22839, 22868, 
    23081, 23484, 24343, 25450, 26945, 22034, 25522, 26323, 25988, 25583, 
    25015, 24508,
  17223, 17416, 22455, 24067, 24933, 24512, 23521, 23074, 22868, 22952, 
    23073, 23560, 24452, 25560, 26594, 22030, 25473, 26257, 25988, 25403, 
    24888, 24382,
  17983, 18102, 22792, 24236, 24991, 24472, 23486, 23063, 22872, 22964, 
    23099, 23538, 24490, 25576, 26703, 22230, 25454, 26338, 25960, 25509, 
    24933, 24429,
  19291, 19330, 23535, 24594, 25042, 24431, 23428, 22983, 22869, 22866, 
    23045, 23576, 24423, 25690, 27040, 22999, 25679, 26273, 25934, 25491, 
    24901, 24389,
  20770, 20760, 24378, 25071, 25177, 24437, 23452, 23054, 22890, 22976, 
    23054, 23604, 24569, 25767, 26645, 24084, 26089, 26295, 25962, 25454, 
    24863, 24276,
  22009, 21988, 24905, 25315, 25206, 24403, 23425, 23019, 22908, 22953, 
    23148, 23579, 24411, 26009, 26766, 24627, 26096, 26301, 25893, 25441, 
    24933, 24243,
  22777, 22752, 25048, 25324, 25111, 24322, 23411, 23005, 22899, 22999, 
    23038, 23508, 24426, 25898, 26982, 24591, 26076, 26360, 26024, 25522, 
    24946, 24450,
  23108, 23066, 25058, 25362, 25123, 24286, 23404, 22967, 22917, 22939, 
    23112, 23658, 24631, 26051, 26389, 24467, 26001, 26288, 25969, 25498, 
    24947, 24497,
  23215, 23151, 25025, 25302, 25121, 24281, 23359, 22982, 22940, 22945, 
    23178, 23735, 24644, 25944, 26953, 24386, 26053, 26281, 25935, 25474, 
    24864, 24397,
  23297, 23230, 25106, 25313, 25058, 24264, 23353, 22956, 22891, 22974, 
    23152, 23722, 24540, 25821, 26944, 24413, 26059, 26246, 25859, 25449, 
    24903, 24304,
  23433, 23385, 25175, 25321, 25032, 24183, 23297, 22982, 22895, 22966, 
    23176, 23646, 24570, 25872, 27228, 24572, 26196, 26159, 25749, 25381, 
    24706, 24271,
  23600, 23588, 25152, 25322, 24998, 24121, 23280, 22962, 22889, 22940, 
    23193, 23768, 24637, 25994, 27218, 24525, 26072, 26051, 25722, 25244, 
    24707, 24238,
  23732, 23748, 25180, 25328, 24935, 24116, 23253, 22977, 22939, 23061, 
    23287, 23786, 24701, 25985, 27216, 24329, 25985, 26029, 25632, 25220, 
    24631, 24125,
  23706, 23704, 25279, 25330, 24913, 24013, 23225, 22972, 22927, 23015, 
    23207, 23637, 24793, 26231, 27264, 24368, 26122, 25943, 25578, 25084, 
    24554, 24045,
  23432, 23332, 25378, 25365, 24850, 23954, 23191, 22986, 22942, 22998, 
    23199, 23787, 24783, 25959, 27035, 24328, 26066, 25957, 25523, 25115, 
    24523, 24052,
  23033, 22796, 25346, 25271, 24793, 23904, 23160, 22958, 22890, 22964, 
    23302, 23843, 24941, 26135, 27170, 24286, 26128, 25959, 25585, 25103, 
    24492, 23939,
  22838, 22535, 25336, 25239, 24699, 23820, 23136, 22919, 22902, 23019, 
    23237, 23855, 24939, 26374, 26882, 24196, 26184, 25929, 25613, 25078, 
    24467, 23940,
  28412, 28313, 27772, 27045, 25747, 24144, 22744, 22225, 22136, 22462, 
    22947, 23620, 24574, 25816, 26888, 28609, 28497, 27271, 26654, 25838, 
    24792, 23869,
  28383, 28297, 27754, 27018, 25826, 24207, 22799, 22231, 22156, 22502, 
    22875, 23590, 24566, 25729, 26674, 28497, 28310, 27041, 26281, 25596, 
    24576, 23789,
  28308, 28262, 27673, 27060, 25912, 24409, 22889, 22319, 22142, 22484, 
    22981, 23549, 24512, 25695, 26562, 28307, 27919, 26694, 26006, 25378, 
    24423, 23655,
  28213, 28215, 27638, 27093, 25949, 24462, 22976, 22348, 22182, 22467, 
    22880, 23538, 24571, 25746, 26723, 28201, 27657, 26385, 25729, 25124, 
    24384, 23635,
  28112, 28131, 27615, 27035, 26015, 24580, 23048, 22359, 22182, 22506, 
    22917, 23573, 24662, 25687, 26868, 28051, 27476, 26232, 25571, 25049, 
    24308, 23655,
  28002, 27980, 27507, 26996, 25998, 24596, 23069, 22477, 22184, 22506, 
    22895, 23560, 24523, 25792, 26635, 27967, 27284, 26168, 25578, 25123, 
    24377, 23827,
  27857, 27765, 27285, 26840, 25951, 24607, 23169, 22462, 22225, 22475, 
    22843, 23538, 24590, 25801, 26921, 27559, 26979, 26088, 25619, 25079, 
    24408, 23734,
  27647, 27513, 27001, 26584, 25837, 24599, 23190, 22523, 22228, 22488, 
    22868, 23504, 24439, 25435, 26607, 26967, 26481, 25872, 25564, 25117, 
    24358, 23807,
  27380, 27249, 26646, 26387, 25728, 24629, 23221, 22550, 22277, 22471, 
    22885, 23514, 24291, 25757, 26732, 26201, 25337, 25346, 25192, 24812, 
    24287, 23740,
  27128, 27005, 26404, 26231, 25746, 24635, 23293, 22585, 22210, 22474, 
    22879, 23499, 24416, 25437, 26660, 25641, 23485, 24480, 24771, 24650, 
    24217, 23706,
  26973, 26843, 26428, 26260, 25757, 24727, 23352, 22617, 22327, 22516, 
    22768, 23471, 24453, 25656, 26598, 25818, 24790, 25107, 25053, 24755, 
    24229, 23752,
  26949, 26825, 26595, 26385, 25834, 24783, 23377, 22623, 22314, 22556, 
    22830, 23551, 24359, 25493, 26865, 26278, 25809, 25540, 25287, 24867, 
    24312, 23618,
  27033, 26951, 26775, 26579, 25974, 24861, 23435, 22669, 22349, 22536, 
    22770, 23389, 24248, 25712, 26450, 26732, 26201, 25684, 25356, 24923, 
    24330, 23718,
  27171, 27138, 26973, 26720, 26117, 24920, 23522, 22693, 22346, 22484, 
    22901, 23439, 24400, 25614, 26457, 27101, 26629, 25900, 25438, 25003, 
    24298, 23825,
  27304, 27288, 27087, 26817, 26137, 24981, 23522, 22760, 22372, 22478, 
    22852, 23421, 24213, 25332, 26588, 27244, 26535, 25732, 25383, 24903, 
    24298, 23798,
  27386, 27354, 27107, 26860, 26148, 25006, 23580, 22778, 22404, 22520, 
    22892, 23396, 24358, 25553, 26604, 27281, 26493, 25726, 25334, 24841, 
    24285, 23757,
  27391, 27346, 27120, 26851, 26207, 25006, 23622, 22810, 22439, 22472, 
    22732, 23352, 24279, 25685, 26864, 27320, 26479, 25754, 25293, 24872, 
    24304, 23804,
  27326, 27291, 27053, 26787, 26199, 25054, 23601, 22833, 22430, 22563, 
    22823, 23444, 24323, 25560, 26828, 27275, 26349, 25668, 25237, 24803, 
    24303, 23823,
  27220, 27199, 27092, 26787, 26240, 25121, 23677, 22883, 22468, 22534, 
    22823, 23357, 24313, 25541, 26449, 27298, 26492, 25747, 25375, 24833, 
    24335, 23816,
  27093, 27072, 27006, 26806, 26248, 25129, 23701, 22883, 22456, 22499, 
    22947, 23420, 24059, 25401, 26495, 27362, 26778, 26035, 25581, 25094, 
    24404, 23889,
  26950, 26916, 26997, 26793, 26256, 25112, 23708, 22912, 22482, 22545, 
    22771, 23448, 24197, 25268, 26599, 27343, 26859, 26187, 25664, 25225, 
    24525, 23836,
  26792, 26755, 26951, 26739, 26173, 25134, 23746, 22950, 22531, 22562, 
    22768, 23311, 24226, 25338, 26553, 27273, 26654, 26135, 25712, 25224, 
    24601, 23902,
  26649, 26628, 26815, 26676, 26193, 25170, 23787, 22941, 22528, 22547, 
    22921, 23358, 24253, 25366, 26759, 27212, 26772, 26279, 25835, 25305, 
    24613, 24002,
  26577, 26577, 26832, 26735, 26250, 25204, 23805, 22947, 22519, 22553, 
    22898, 23368, 24295, 25396, 26494, 27288, 27039, 26388, 25904, 25268, 
    24645, 23955,
  26617, 26621, 26901, 26739, 26313, 25235, 23846, 23000, 22519, 22541, 
    22847, 23393, 24312, 25270, 26475, 27424, 27076, 26359, 25863, 25224, 
    24600, 24008,
  26755, 26744, 26951, 26822, 26310, 25277, 23863, 23005, 22568, 22564, 
    22844, 23368, 24152, 25293, 26907, 27410, 27107, 26395, 25960, 25379, 
    24702, 24041,
  26924, 26893, 27089, 26826, 26229, 25237, 23856, 23020, 22592, 22555, 
    22877, 23254, 24257, 25233, 26492, 27324, 27001, 26373, 25966, 25435, 
    24657, 24067,
  27042, 26992, 27063, 26822, 26232, 25251, 23925, 23046, 22618, 22549, 
    22792, 23291, 24250, 25512, 26647, 27321, 26851, 26395, 26042, 25559, 
    24771, 24061,
  27046, 26977, 27096, 26876, 26279, 25237, 23939, 23052, 22597, 22546, 
    22926, 23342, 24119, 25251, 26460, 27413, 27188, 26590, 26090, 25559, 
    24841, 24134,
  26914, 26831, 27071, 26862, 26301, 25293, 23925, 23040, 22600, 22528, 
    22823, 23286, 24323, 25384, 26341, 27478, 27325, 26654, 26256, 25701, 
    24930, 24301,
  26678, 26598, 26949, 26757, 26329, 25296, 23939, 23093, 22661, 22560, 
    22877, 23316, 24220, 25333, 26110, 27400, 27307, 26719, 26310, 25764, 
    25031, 24307,
  26407, 26340, 26850, 26684, 26229, 25265, 23939, 23111, 22617, 22574, 
    22859, 23346, 24289, 25216, 26540, 27274, 27251, 26704, 26290, 25844, 
    25108, 24407,
  26149, 26083, 26644, 26568, 26207, 25253, 23994, 23128, 22699, 22640, 
    22811, 23323, 24135, 25171, 26399, 27169, 27089, 26589, 26269, 25819, 
    25184, 24534,
  25896, 25824, 26560, 26498, 26151, 25245, 23966, 23131, 22676, 22639, 
    22868, 23346, 24128, 25400, 26585, 27049, 27001, 26632, 26262, 25838, 
    25235, 24568,
  25625, 25564, 26497, 26407, 26089, 25248, 23942, 23148, 22675, 22622, 
    22856, 23382, 24175, 25416, 26322, 26920, 26926, 26582, 26235, 25782, 
    25260, 24607,
  25358, 25329, 26249, 26304, 26026, 25234, 23987, 23169, 22701, 22590, 
    22785, 23323, 24086, 25427, 26426, 26809, 26876, 26509, 26172, 25775, 
    25228, 24620,
  25158, 25148, 26114, 26185, 26017, 25214, 23959, 23160, 22690, 22573, 
    22807, 23315, 24212, 25392, 26064, 26628, 26782, 26422, 26213, 25800, 
    25273, 24647,
  25071, 25039, 25873, 26101, 25975, 25152, 23969, 23151, 22727, 22630, 
    22745, 23371, 24051, 25327, 26760, 26426, 26571, 26322, 25999, 25676, 
    25094, 24660,
  25078, 24994, 25904, 26088, 25917, 25183, 23955, 23172, 22692, 22622, 
    22813, 23231, 24139, 25357, 26054, 26285, 26503, 26220, 25896, 25570, 
    25120, 24701,
  25102, 24981, 26091, 26175, 25966, 25197, 24035, 23186, 22698, 22641, 
    22807, 23363, 24085, 25409, 26190, 26269, 26553, 26249, 25944, 25632, 
    25164, 24634,
  25074, 24962, 26038, 26207, 26014, 25239, 24001, 23221, 22715, 22624, 
    22881, 23333, 24147, 25283, 26578, 26207, 26503, 26090, 25847, 25501, 
    25087, 24580,
  25008, 24940, 25957, 26164, 26038, 25228, 23993, 23186, 22765, 22638, 
    22884, 23404, 24124, 25245, 26226, 26038, 26596, 26249, 25903, 25563, 
    25043, 24613,
  24998, 24975, 25893, 26113, 26040, 25214, 23972, 23186, 22733, 22667, 
    22864, 23307, 24152, 25190, 26518, 25885, 26682, 26271, 25929, 25563, 
    25176, 24714,
  25127, 25126, 25995, 26175, 26079, 25275, 24018, 23186, 22791, 22613, 
    22852, 23261, 24258, 25264, 26299, 25974, 26682, 26285, 25901, 25482, 
    25017, 24673,
  25374, 25369, 26190, 26323, 26106, 25312, 23997, 23192, 22733, 22589, 
    22855, 23279, 24285, 25546, 26479, 26110, 26826, 26357, 25978, 25507, 
    25042, 24546,
  25622, 25603, 26354, 26447, 26189, 25259, 24007, 23212, 22748, 22650, 
    22875, 23239, 24206, 25320, 26457, 26242, 26807, 26307, 25937, 25489, 
    24992, 24479,
  25750, 25736, 26537, 26541, 26169, 25281, 23959, 23254, 22765, 22630, 
    22938, 23296, 24186, 25310, 26032, 26422, 26764, 26226, 25804, 25352, 
    24852, 24446,
  25721, 25750, 26504, 26525, 26189, 25233, 24011, 23221, 22762, 22655, 
    22904, 23317, 24085, 25164, 26190, 26431, 26632, 26176, 25716, 25320, 
    24782, 24379,
  25603, 25689, 26456, 26528, 26212, 25273, 24049, 23242, 22756, 22664, 
    22869, 23332, 24265, 25271, 26539, 26375, 26789, 26249, 25743, 25345, 
    24820, 24472,
  25506, 25610, 26375, 26450, 26129, 25320, 24000, 23242, 22806, 22699, 
    22955, 23312, 24110, 25204, 26464, 26229, 26851, 26393, 25881, 25432, 
    24750, 24286,
  25492, 25559, 26266, 26342, 26146, 25255, 23996, 23274, 22754, 22661, 
    22964, 23269, 24243, 25366, 26294, 26122, 26751, 26415, 25916, 25370, 
    24756, 24339,
  25528, 25543, 26253, 26401, 26135, 25281, 24025, 23251, 22803, 22721, 
    22964, 23332, 24036, 25254, 26420, 26088, 26653, 26401, 25806, 25308, 
    24731, 24259,
  25513, 25520, 26360, 26420, 26146, 25236, 24000, 23221, 22771, 22741, 
    22912, 23378, 24050, 25481, 26134, 26213, 26721, 26285, 25840, 25333, 
    24705, 24179,
  25358, 25414, 26385, 26422, 26112, 25228, 23972, 23266, 22818, 22748, 
    22952, 23337, 24083, 25204, 26139, 26291, 26889, 26328, 25799, 25333, 
    24731, 24118,
  25052, 25168, 26142, 26312, 26072, 25256, 23969, 23245, 22844, 22696, 
    22947, 23449, 24011, 25071, 26585, 26049, 26901, 26451, 25937, 25364, 
    24750, 24172,
  24629, 24770, 25954, 26157, 25992, 25219, 23979, 23233, 22800, 22667, 
    22896, 23381, 24280, 25238, 26757, 25692, 26671, 26567, 26129, 25495, 
    24769, 24192,
  24095, 24216, 25612, 25910, 25929, 25166, 23990, 23195, 22865, 22699, 
    22913, 23381, 24260, 25430, 26409, 25403, 26876, 26704, 26144, 25532, 
    24807, 24166,
  23377, 23482, 25193, 25685, 25831, 25172, 23973, 23245, 22816, 22736, 
    22913, 23384, 24194, 25357, 26554, 25104, 26757, 26732, 26185, 25620, 
    24826, 24239,
  22394, 22538, 24960, 25499, 25704, 25090, 23997, 23207, 22821, 22696, 
    22938, 23333, 24162, 25274, 26438, 24781, 26540, 26726, 26254, 25707, 
    24967, 24333,
  21177, 21421, 24737, 25394, 25657, 25099, 23921, 23195, 22822, 22733, 
    22853, 23371, 24256, 25497, 26462, 24608, 26466, 26820, 26351, 25738, 
    25088, 24373,
  19941, 20293, 23964, 24880, 25453, 25046, 23917, 23204, 22830, 22791, 
    22939, 23463, 24226, 25472, 26278, 23753, 26142, 26748, 26331, 25806, 
    25012, 24427,
  19010, 19428, 22904, 24193, 25142, 24928, 23935, 23204, 22839, 22751, 
    22976, 23394, 24128, 25432, 26484, 22361, 25028, 26473, 26304, 25775, 
    25063, 24407,
  18643, 19072, 22770, 24134, 25107, 24931, 23869, 23213, 22801, 22725, 
    23028, 23338, 24291, 25444, 26448, 22294, 25177, 26553, 26357, 25906, 
    25120, 24447,
  18891, 19281, 23069, 24315, 25133, 24903, 23866, 23202, 22828, 22780, 
    23028, 23488, 24227, 25477, 26795, 22764, 25420, 26582, 26345, 25925, 
    25177, 24514,
  19568, 19876, 23396, 24436, 25196, 24881, 23845, 23146, 22866, 22777, 
    23005, 23425, 24375, 25383, 26470, 23011, 25427, 26531, 26345, 25900, 
    25254, 24588,
  20369, 20580, 23845, 24759, 25316, 24892, 23859, 23167, 22860, 22818, 
    23028, 23367, 24200, 25333, 26970, 23557, 25582, 26597, 26351, 25944, 
    25229, 24608,
  21035, 21189, 24271, 24991, 25382, 24872, 23804, 23158, 22899, 22778, 
    22937, 23425, 24313, 25300, 26489, 24033, 25856, 26560, 26351, 25901, 
    25204, 24602,
  21466, 21626, 24312, 24977, 25377, 24839, 23786, 23152, 22817, 22729, 
    23068, 23451, 24198, 25381, 26523, 24055, 25862, 26582, 26318, 25882, 
    25159, 24669,
  21705, 21893, 24236, 24918, 25340, 24817, 23790, 23141, 22823, 22801, 
    22940, 23431, 24144, 25417, 26747, 23932, 25707, 26532, 26221, 25801, 
    25172, 24636,
  21836, 22013, 24246, 24967, 25283, 24845, 23786, 23182, 22820, 22807, 
    23080, 23393, 24304, 25507, 26672, 23957, 25713, 26496, 26215, 25696, 
    25032, 24442,
  21900, 22024, 24449, 25069, 25325, 24814, 23717, 23123, 22838, 22793, 
    22975, 23398, 24262, 25296, 26625, 24040, 25676, 26467, 26118, 25726, 
    25077, 24496,
  21889, 21978, 24490, 25147, 25329, 24775, 23707, 23132, 22885, 22787, 
    22995, 23431, 24262, 25405, 26456, 24196, 25664, 26460, 26194, 25659, 
    25007, 24449,
  21791, 21904, 24411, 25112, 25303, 24739, 23704, 23141, 22862, 22908, 
    23006, 23442, 24322, 25375, 26616, 24224, 25869, 26475, 26119, 25628, 
    25065, 24609,
  21598, 21773, 24340, 25048, 25295, 24728, 23714, 23133, 22873, 22865, 
    22987, 23462, 24359, 25660, 26632, 24254, 25994, 26446, 26070, 25690, 
    25039, 24570,
  21282, 21513, 24269, 24975, 25278, 24672, 23645, 23089, 22859, 22851, 
    23036, 23432, 24263, 25706, 26599, 24164, 26013, 26482, 26112, 25715, 
    25084, 24550,
  20799, 21055, 24107, 24941, 25203, 24683, 23631, 23089, 22865, 22906, 
    23116, 23435, 24401, 25454, 26771, 23983, 25820, 26439, 26153, 25716, 
    25193, 24677,
  20122, 20379, 23859, 24774, 25135, 24596, 23631, 23083, 22912, 22797, 
    23076, 23481, 24476, 25662, 26803, 23650, 25771, 26432, 26147, 25759, 
    25187, 24798,
  19286, 19539, 23299, 24470, 25075, 24585, 23611, 23107, 22863, 22984, 
    23062, 23471, 24363, 25716, 26757, 23107, 25659, 26338, 26113, 25691, 
    25136, 24718,
  18445, 18695, 22770, 24231, 24998, 24572, 23559, 23054, 22851, 22912, 
    22985, 23491, 24471, 25595, 26726, 22392, 25429, 26367, 26078, 25635, 
    25111, 24684,
  17869, 18101, 22474, 24078, 24912, 24502, 23566, 23075, 22857, 22884, 
    23037, 23563, 24447, 25651, 26794, 22033, 25367, 26317, 26024, 25679, 
    25067, 24525,
  17842, 18013, 22563, 24137, 24918, 24552, 23573, 23067, 22869, 22875, 
    23017, 23565, 24378, 25714, 26445, 21976, 25311, 26303, 25969, 25555, 
    24851, 24291,
  18479, 18554, 22756, 24250, 24921, 24477, 23539, 23041, 22881, 22954, 
    23080, 23599, 24502, 25637, 26585, 22098, 25429, 26346, 26010, 25518, 
    24883, 24385,
  19633, 19618, 23394, 24549, 25050, 24412, 23480, 23032, 22920, 22960, 
    23157, 23644, 24482, 25619, 26721, 22817, 25579, 26310, 25962, 25550, 
    24985, 24412,
  20957, 20895, 24289, 24998, 25122, 24435, 23526, 23038, 22894, 22954, 
    23118, 23637, 24408, 25801, 26660, 23854, 25915, 26304, 26024, 25612, 
    25017, 24479,
  22079, 22013, 24892, 25268, 25219, 24371, 23467, 23017, 22923, 22954, 
    23104, 23640, 24529, 25588, 26656, 24495, 26082, 26304, 26066, 25631, 
    25093, 24600,
  22792, 22728, 25034, 25349, 25165, 24374, 23435, 23018, 22873, 22948, 
    23124, 23666, 24352, 25932, 26756, 24601, 26120, 26318, 25997, 25693, 
    25126, 24587,
  23119, 23045, 25004, 25354, 25202, 24337, 23391, 23015, 22924, 22961, 
    23061, 23674, 24384, 25854, 26998, 24517, 26021, 26310, 25997, 25613, 
    25120, 24687,
  23238, 23154, 25123, 25359, 25105, 24288, 23377, 22992, 22912, 22958, 
    23164, 23555, 24565, 25647, 26876, 24466, 26096, 26275, 26039, 25607, 
    25177, 24587,
  23323, 23246, 25098, 25362, 25085, 24195, 23343, 23021, 22927, 22978, 
    23094, 23659, 24621, 26050, 26984, 24477, 26139, 26260, 25895, 25520, 
    25031, 24527,
  23457, 23393, 25129, 25370, 25051, 24184, 23353, 23004, 22945, 22990, 
    23156, 23750, 24784, 25920, 26928, 24476, 26132, 26160, 25874, 25514, 
    24898, 24414,
  23642, 23592, 25172, 25422, 25008, 24109, 23319, 23004, 22951, 23033, 
    23222, 23748, 24573, 26157, 26882, 24484, 26090, 26110, 25757, 25471, 
    24867, 24355,
  23824, 23787, 25316, 25352, 24954, 24089, 23253, 22978, 22922, 22976, 
    23168, 23723, 24679, 25785, 27110, 24397, 26078, 26074, 25701, 25279, 
    24651, 24255,
  23874, 23827, 25352, 25379, 24917, 24014, 23198, 22979, 22948, 22974, 
    23348, 23781, 24679, 25960, 26946, 24539, 26071, 26010, 25578, 25130, 
    24588, 24142,
  23680, 23562, 25426, 25396, 24886, 23978, 23205, 23014, 22955, 22971, 
    23254, 23777, 24724, 26022, 27098, 24553, 26122, 25916, 25517, 25074, 
    24550, 24102,
  23341, 23114, 25395, 25320, 24792, 23869, 23153, 22985, 22958, 23014, 
    23226, 23891, 24800, 26057, 27045, 24491, 26090, 25859, 25469, 25099, 
    24525, 23942,
  23168, 22885, 25438, 25329, 24715, 23807, 23112, 22953, 22935, 22992, 
    23291, 23846, 24877, 26054, 27234, 24374, 26072, 25881, 25490, 25056, 
    24424, 23963,
  28331, 28186, 27732, 26990, 25728, 24126, 22746, 22245, 22110, 22479, 
    23041, 23608, 24653, 25660, 26709, 28507, 28128, 26876, 26266, 25514, 
    24482, 23668,
  28292, 28158, 27665, 26987, 25807, 24230, 22808, 22268, 22162, 22567, 
    22927, 23499, 24554, 25609, 26615, 28335, 27891, 26573, 26004, 25303, 
    24444, 23707,
  28199, 28099, 27574, 26942, 25854, 24322, 22933, 22323, 22194, 22547, 
    22927, 23569, 24611, 25976, 26706, 28141, 27549, 26328, 25742, 25135, 
    24298, 23580,
  28094, 28043, 27500, 26947, 25899, 24429, 22975, 22362, 22223, 22463, 
    22935, 23554, 24337, 25622, 26939, 27984, 27306, 26069, 25467, 24862, 
    24234, 23546,
  27997, 27970, 27484, 26922, 25962, 24504, 23058, 22423, 22188, 22529, 
    22963, 23559, 24303, 25703, 26549, 27897, 27313, 26126, 25543, 24948, 
    24246, 23539,
  27898, 27841, 27439, 26885, 25962, 24523, 23068, 22423, 22211, 22472, 
    22849, 23500, 24393, 25606, 26803, 27763, 27256, 26184, 25679, 25004, 
    24290, 23659,
  27766, 27651, 27173, 26723, 25862, 24574, 23179, 22446, 22257, 22474, 
    22800, 23500, 24405, 25570, 26839, 27364, 26896, 26054, 25618, 25028, 
    24347, 23705,
  27575, 27432, 26889, 26446, 25790, 24601, 23157, 22473, 22231, 22497, 
    22840, 23606, 24474, 25370, 26381, 26621, 26254, 25823, 25452, 25034, 
    24397, 23825,
  27333, 27212, 26562, 26346, 25690, 24587, 23244, 22572, 22245, 22516, 
    22800, 23489, 24472, 25579, 27014, 25957, 24762, 25138, 25129, 24786, 
    24257, 23812,
  27104, 27015, 26485, 26260, 25698, 24676, 23310, 22611, 22257, 22476, 
    22939, 23520, 24543, 25533, 26519, 25824, 23911, 24763, 24901, 24773, 
    24314, 23745,
  26959, 26877, 26531, 26338, 25787, 24730, 23368, 22584, 22274, 22524, 
    22882, 23506, 24572, 25493, 26285, 26156, 25166, 25282, 25114, 24884, 
    24289, 23791,
  26933, 26846, 26647, 26443, 25870, 24760, 23393, 22648, 22323, 22432, 
    22867, 23390, 24382, 25523, 26167, 26541, 25595, 25461, 25238, 24859, 
    24313, 23777,
  27003, 26930, 26817, 26582, 25984, 24881, 23452, 22674, 22352, 22506, 
    22850, 23476, 24409, 25516, 26521, 26807, 26074, 25606, 25313, 24934, 
    24288, 23837,
  27124, 27080, 26959, 26657, 26084, 24903, 23479, 22701, 22366, 22481, 
    22850, 23514, 24478, 25497, 26790, 27104, 26714, 25929, 25464, 24952, 
    24408, 23890,
  27254, 27219, 27089, 26790, 26104, 25006, 23527, 22748, 22396, 22532, 
    22830, 23445, 24278, 25537, 26722, 27273, 26876, 26117, 25574, 25038, 
    24395, 23830,
  27353, 27297, 27114, 26819, 26132, 24978, 23586, 22783, 22380, 22517, 
    22829, 23442, 24265, 25420, 26382, 27312, 26626, 25806, 25436, 24877, 
    24274, 23803,
  27387, 27311, 27144, 26806, 26184, 25065, 23631, 22821, 22462, 22517, 
    22826, 23358, 24258, 25436, 26510, 27290, 26248, 25525, 25195, 24777, 
    24254, 23762,
  27341, 27275, 27060, 26810, 26190, 24989, 23638, 22824, 22468, 22485, 
    22860, 23467, 24265, 25343, 26438, 27243, 26328, 25547, 25222, 24845, 
    24299, 23829,
  27224, 27189, 27026, 26846, 26198, 25101, 23679, 22864, 22447, 22516, 
    22834, 23444, 24304, 25352, 26367, 27265, 26596, 25799, 25374, 24975, 
    24298, 23808,
  27058, 27045, 27020, 26784, 26181, 25106, 23672, 22861, 22470, 22504, 
    22851, 23352, 24297, 25478, 26476, 27326, 26894, 26072, 25560, 25124, 
    24463, 23908,
  26861, 26846, 26984, 26741, 26172, 25126, 23720, 22902, 22514, 22516, 
    22794, 23362, 24296, 25403, 26476, 27301, 26826, 26209, 25746, 25292, 
    24539, 24002,
  26656, 26629, 26857, 26635, 26140, 25075, 23769, 22923, 22560, 22521, 
    22776, 23519, 24308, 25682, 26582, 27115, 26521, 26129, 25773, 25291, 
    24590, 24068,
  26482, 26456, 26809, 26635, 26151, 25162, 23769, 22937, 22586, 22544, 
    22799, 23346, 24291, 25522, 26485, 27009, 26346, 26115, 25800, 25335, 
    24603, 23934,
  26393, 26377, 26720, 26635, 26179, 25224, 23848, 22996, 22574, 22518, 
    22824, 23455, 24293, 25336, 26510, 27115, 26688, 26259, 25862, 25309, 
    24628, 23987,
  26421, 26403, 26847, 26729, 26251, 25210, 23838, 22978, 22586, 22589, 
    22841, 23376, 24244, 25296, 26595, 27294, 27006, 26447, 25944, 25452, 
    24704, 24060,
  26545, 26506, 26938, 26762, 26220, 25223, 23855, 23022, 22586, 22560, 
    22941, 23452, 24155, 25246, 26318, 27266, 26975, 26418, 25957, 25539, 
    24768, 24141,
  26698, 26635, 26948, 26732, 26223, 25218, 23872, 23069, 22574, 22534, 
    22852, 23335, 24157, 25388, 26622, 27219, 26850, 26432, 26082, 25532, 
    24786, 24154,
  26807, 26730, 26935, 26762, 26263, 25215, 23851, 23054, 22603, 22566, 
    22892, 23378, 24177, 25349, 26544, 27199, 26863, 26439, 26026, 25582, 
    24875, 24193,
  26822, 26734, 26999, 26794, 26274, 25226, 23900, 23054, 22562, 22606, 
    22880, 23373, 24297, 25193, 26497, 27275, 27154, 26569, 26103, 25600, 
    24951, 24273,
  26733, 26632, 27007, 26800, 26323, 25307, 23907, 23063, 22626, 22614, 
    22794, 23291, 24193, 25342, 26551, 27306, 27229, 26604, 26206, 25706, 
    25002, 24447,
  26576, 26467, 26768, 26718, 26207, 25234, 23931, 23110, 22658, 22542, 
    22846, 23408, 24198, 25286, 26553, 27269, 27273, 26699, 26282, 25887, 
    25117, 24534,
  26411, 26299, 26682, 26626, 26240, 25245, 23945, 23095, 22658, 22590, 
    22837, 23286, 24075, 25265, 26307, 27119, 27235, 26641, 26301, 25885, 
    25167, 24514,
  26261, 26151, 26656, 26619, 26191, 25268, 23938, 23127, 22660, 22602, 
    22794, 23425, 24211, 25346, 26274, 27041, 27149, 26663, 26247, 25829, 
    25224, 24534,
  26096, 25997, 26621, 26526, 26168, 25253, 23927, 23156, 22687, 22562, 
    22834, 23309, 24176, 25216, 26582, 26926, 26949, 26590, 26212, 25818, 
    25218, 24594,
  25887, 25814, 26387, 26447, 26119, 25236, 23958, 23156, 22701, 22564, 
    22968, 23392, 24264, 25260, 26376, 26829, 26985, 26554, 26171, 25829, 
    25218, 24661,
  25655, 25614, 26282, 26357, 26104, 25265, 23948, 23177, 22681, 22662, 
    22876, 23311, 24289, 25434, 26269, 26679, 26849, 26453, 26101, 25817, 
    25249, 24727,
  25467, 25436, 26088, 26242, 26034, 25236, 23968, 23197, 22774, 22619, 
    22876, 23369, 24279, 25281, 26616, 26456, 26837, 26409, 26088, 25754, 
    25325, 24707,
  25372, 25319, 25869, 26099, 25950, 25192, 23948, 23197, 22721, 22638, 
    22822, 23420, 24158, 25397, 26766, 26169, 26706, 26301, 25976, 25704, 
    25236, 24714,
  25364, 25275, 25966, 26120, 25965, 25200, 23989, 23206, 22739, 22658, 
    22773, 23341, 24239, 25194, 26810, 26088, 26532, 26250, 25991, 25717, 
    25300, 24754,
  25386, 25281, 26079, 26257, 26001, 25203, 23985, 23171, 22727, 22613, 
    22876, 23318, 24081, 25166, 26118, 26181, 26506, 26243, 25895, 25593, 
    25236, 24774,
  25383, 25300, 26138, 26271, 26032, 25197, 23926, 23176, 22704, 22586, 
    22878, 23381, 24094, 25199, 26422, 26182, 26619, 26250, 25907, 25618, 
    25249, 24928,
  25367, 25325, 26014, 26206, 26067, 25228, 23982, 23173, 22756, 22627, 
    22847, 23366, 24111, 25241, 26570, 26022, 26762, 26351, 25957, 25673, 
    25325, 24928,
  25415, 25410, 25768, 26131, 26004, 25278, 23975, 23247, 22735, 22610, 
    22927, 23340, 24150, 25241, 26313, 25749, 26575, 26344, 25998, 25660, 
    25236, 24854,
  25585, 25596, 25979, 26257, 26099, 25323, 23971, 23185, 22750, 22641, 
    22844, 23272, 24079, 25522, 26494, 25829, 26600, 26322, 25894, 25593, 
    25134, 24780,
  25828, 25840, 26371, 26460, 26188, 25314, 24024, 23191, 22780, 22735, 
    22770, 23350, 24197, 25310, 26421, 26242, 26879, 26387, 25956, 25555, 
    25198, 24746,
  26022, 26031, 26740, 26662, 26276, 25284, 23929, 23200, 22762, 22684, 
    22847, 23274, 24145, 25348, 26506, 26651, 26949, 26344, 25825, 25462, 
    25064, 24593,
  26072, 26092, 26757, 26654, 26229, 25295, 23999, 23241, 22774, 22663, 
    22890, 23310, 24194, 25308, 26269, 26751, 26818, 26221, 25756, 25363, 
    24936, 24465,
  25987, 26040, 26598, 26604, 26222, 25273, 23982, 23197, 22785, 22669, 
    22935, 23345, 24187, 25015, 26356, 26601, 26849, 26300, 25756, 25313, 
    24758, 24459,
  25858, 25952, 26517, 26497, 26196, 25273, 23995, 23217, 22753, 22715, 
    22910, 23421, 24177, 25264, 26720, 26498, 26885, 26300, 25839, 25313, 
    24726, 24305,
  25790, 25897, 26488, 26514, 26213, 25286, 23995, 23253, 22785, 22690, 
    22918, 23345, 24170, 25443, 26378, 26515, 26854, 26307, 25763, 25170, 
    24733, 24225,
  25821, 25903, 26537, 26540, 26210, 25314, 23978, 23208, 22782, 22675, 
    22918, 23325, 24145, 25371, 26492, 26524, 26806, 26228, 25770, 25244, 
    24694, 24285,
  25898, 25953, 26539, 26572, 26245, 25298, 23995, 23253, 22809, 22695, 
    22910, 23264, 24061, 25376, 26448, 26546, 26787, 26228, 25749, 25182, 
    24631, 24238,
  25915, 25987, 26559, 26540, 26159, 25259, 23964, 23217, 22765, 22595, 
    22853, 23300, 24234, 25406, 26401, 26588, 26917, 26337, 25866, 25226, 
    24669, 24238,
  25794, 25919, 26534, 26504, 26128, 25253, 23975, 23232, 22780, 22730, 
    22890, 23401, 24148, 25171, 26625, 26573, 27017, 26488, 25970, 25406, 
    24778, 24251,
  25513, 25676, 26420, 26454, 26122, 25214, 23958, 23217, 22785, 22684, 
    22935, 23356, 24185, 25285, 26360, 26493, 27079, 26553, 26067, 25431, 
    24739, 24191,
  25076, 25230, 26243, 26295, 26065, 25194, 23985, 23268, 22827, 22701, 
    22970, 23392, 24261, 25248, 26460, 26267, 27079, 26662, 26156, 25556, 
    24809, 24218,
  24466, 24583, 25900, 26107, 25985, 25225, 23930, 23212, 22806, 22730, 
    23007, 23404, 24146, 25311, 26550, 25879, 26954, 26698, 26135, 25599, 
    24924, 24278,
  23639, 23744, 25347, 25781, 25876, 25211, 23968, 23206, 22844, 22699, 
    22919, 23419, 24163, 25406, 26535, 25228, 26582, 26698, 26225, 25674, 
    24962, 24352,
  22576, 22736, 24905, 25541, 25729, 25133, 23951, 23215, 22824, 22722, 
    22902, 23397, 24311, 25334, 26300, 24651, 26257, 26726, 26350, 25848, 
    25052, 24486,
  21368, 21629, 24530, 25320, 25679, 25049, 23916, 23206, 22850, 22759, 
    22996, 23384, 24252, 25308, 26422, 24528, 26500, 26799, 26371, 25854, 
    25141, 24593,
  20237, 20594, 23851, 24884, 25415, 25034, 23906, 23197, 22798, 22779, 
    22996, 23405, 24069, 25474, 27026, 23740, 26065, 26676, 26323, 25892, 
    25077, 24486,
  19468, 19873, 23050, 24276, 25163, 24945, 23899, 23198, 22824, 22728, 
    23033, 23534, 24276, 25374, 26475, 22570, 25087, 26503, 26232, 25879, 
    25179, 24533,
  19259, 19657, 23085, 24335, 25155, 24905, 23843, 23204, 22860, 22765, 
    22919, 23326, 24272, 25344, 26232, 22695, 25405, 26575, 26295, 25879, 
    25135, 24547,
  19597, 19945, 23453, 24556, 25218, 24878, 23850, 23212, 22848, 22797, 
    22996, 23428, 24354, 25381, 26310, 23151, 25642, 26576, 26357, 25867, 
    25199, 24634,
  20266, 20531, 23839, 24699, 25278, 24897, 23879, 23213, 22883, 22786, 
    23034, 23509, 24316, 25241, 26760, 23408, 25529, 26560, 26329, 25954, 
    25263, 24681,
  20967, 21152, 24257, 24963, 25381, 24897, 23816, 23154, 22828, 22800, 
    22966, 23405, 24257, 25405, 26500, 23975, 25891, 26619, 26460, 25948, 
    25314, 24748,
  21493, 21643, 24382, 25057, 25418, 24900, 23840, 23136, 22851, 22783, 
    23034, 23398, 24354, 25488, 26468, 24240, 25997, 26598, 26392, 25954, 
    25193, 24702,
  21800, 21964, 24313, 25087, 25347, 24892, 23806, 23136, 22840, 22824, 
    23111, 23484, 24310, 25676, 26867, 24145, 25866, 26569, 26310, 25899, 
    25187, 24655,
  21958, 22136, 24240, 25012, 25356, 24825, 23789, 23140, 22872, 22844, 
    22969, 23495, 24228, 25460, 26809, 24017, 25779, 26562, 26268, 25763, 
    25143, 24629,
  22035, 22183, 24288, 25036, 25361, 24817, 23734, 23146, 22878, 22821, 
    22997, 23465, 24362, 25338, 26485, 24016, 25692, 26454, 26137, 25719, 
    25111, 24562,
  22045, 22140, 24519, 25179, 25350, 24811, 23744, 23152, 22861, 22913, 
    23029, 23561, 24140, 25514, 26459, 24281, 25854, 26490, 26241, 25719, 
    25162, 24662,
  21974, 22054, 24598, 25206, 25384, 24795, 23737, 23143, 22885, 22813, 
    23029, 23473, 24239, 25514, 26673, 24506, 26029, 26510, 26207, 25713, 
    25207, 24696,
  21837, 21961, 24502, 25157, 25339, 24752, 23678, 23120, 22841, 22865, 
    23129, 23544, 24293, 25454, 26629, 24486, 26228, 26534, 26214, 25769, 
    25207, 24736,
  21664, 21854, 24263, 25026, 25259, 24747, 23724, 23103, 22882, 22851, 
    23118, 23445, 24278, 25596, 27044, 24307, 26085, 26497, 26200, 25807, 
    25284, 24770,
  21452, 21689, 24286, 25002, 25259, 24705, 23661, 23100, 22876, 22882, 
    23010, 23519, 24261, 25522, 26595, 24218, 26066, 26482, 26131, 25764, 
    25208, 24710,
  21143, 21406, 24324, 25018, 25213, 24652, 23647, 23073, 22862, 22897, 
    23042, 23476, 24378, 25635, 26916, 24240, 26066, 26469, 26145, 25795, 
    25182, 24750,
  20664, 20949, 24243, 24986, 25239, 24652, 23617, 23106, 22901, 22871, 
    23105, 23491, 24481, 25645, 26615, 24092, 26017, 26368, 26118, 25664, 
    25138, 24570,
  20007, 20310, 23836, 24782, 25125, 24669, 23613, 23150, 22871, 22886, 
    23168, 23497, 24519, 25599, 26510, 23598, 25893, 26412, 26070, 25701, 
    25126, 24684,
  19292, 19590, 23192, 24459, 25071, 24599, 23617, 23074, 22930, 22909, 
    23100, 23575, 24270, 25541, 26685, 22870, 25551, 26382, 26139, 25721, 
    25215, 24671,
  18765, 19016, 22924, 24314, 25025, 24557, 23558, 23057, 22913, 22909, 
    23111, 23622, 24349, 25448, 26401, 22365, 25395, 26268, 26029, 25665, 
    24993, 24471,
  18688, 18847, 22946, 24338, 24968, 24527, 23513, 23089, 22899, 22872, 
    23109, 23548, 24293, 25701, 26763, 22253, 25389, 26260, 25967, 25541, 
    24993, 24417,
  19177, 19225, 23026, 24371, 25011, 24460, 23524, 23060, 22861, 22930, 
    23074, 23584, 24460, 25567, 26417, 22199, 25265, 26282, 25967, 25461, 
    24936, 24391,
  20117, 20076, 23525, 24637, 25020, 24427, 23517, 23069, 22902, 22956, 
    23140, 23551, 24456, 25744, 26457, 22648, 25352, 26376, 25995, 25597, 
    25000, 24485,
  21216, 21139, 24235, 24976, 25080, 24387, 23455, 23067, 22914, 22950, 
    23140, 23694, 24587, 25856, 26693, 23567, 25676, 26282, 26023, 25654, 
    25076, 24539,
  22168, 22095, 24812, 25259, 25189, 24430, 23424, 23040, 22888, 22968, 
    23089, 23590, 24528, 25629, 26660, 24342, 26068, 26341, 26051, 25728, 
    25159, 24566,
  22795, 22732, 24988, 25345, 25169, 24379, 23424, 23052, 22920, 22974, 
    23124, 23588, 24560, 25558, 27032, 24537, 26168, 26304, 25989, 25710, 
    25192, 24653,
  23109, 23047, 25076, 25375, 25112, 24340, 23424, 23050, 22929, 22986, 
    23221, 23714, 24580, 25940, 26956, 24481, 26104, 26313, 26010, 25629, 
    25109, 24647,
  23250, 23190, 25109, 25386, 25121, 24301, 23387, 23038, 22935, 23009, 
    23204, 23745, 24674, 25682, 27075, 24458, 26149, 26254, 25982, 25556, 
    25001, 24513,
  23360, 23306, 25112, 25394, 25101, 24248, 23352, 23018, 22918, 23009, 
    23267, 23700, 24795, 25803, 27249, 24430, 26154, 26154, 25865, 25550, 
    24969, 24427,
  23514, 23451, 25231, 25375, 25046, 24201, 23345, 23045, 22924, 23018, 
    23171, 23698, 24743, 25735, 27176, 24491, 26056, 26126, 25825, 25426, 
    24830, 24333,
  23726, 23642, 25285, 25383, 25032, 24156, 23290, 23027, 22971, 23027, 
    23197, 23784, 24647, 26187, 26960, 24507, 26125, 26104, 25797, 25401, 
    24850, 24320,
  23947, 23856, 25341, 25378, 24970, 24084, 23259, 23034, 22969, 23004, 
    23234, 23767, 24776, 25894, 27174, 24471, 26112, 26090, 25735, 25370, 
    24729, 24200,
  24044, 23956, 25480, 25394, 24913, 24044, 23249, 23040, 22939, 22999, 
    23208, 23828, 24722, 26207, 27001, 24604, 26162, 26004, 25639, 25215, 
    24590, 24194,
  23891, 23773, 25445, 25386, 24853, 23963, 23246, 22996, 22975, 23016, 
    23226, 23752, 24971, 26104, 26920, 24665, 26150, 25910, 25522, 25061, 
    24507, 24041,
  23583, 23395, 25447, 25355, 24802, 23896, 23170, 22984, 23019, 23108, 
    23294, 23752, 24907, 26346, 27154, 24670, 26175, 25910, 25461, 25042, 
    24527, 24021,
  23421, 23194, 25372, 25311, 24764, 23835, 23197, 22949, 22967, 23063, 
    23318, 23788, 24860, 25990, 27284, 24559, 26138, 25817, 25399, 24894, 
    24375, 23881,
  28234, 28081, 27593, 26910, 25707, 24155, 22772, 22285, 22142, 22524, 
    22934, 23603, 24616, 25901, 26572, 28297, 27720, 26607, 25982, 25281, 
    24308, 23626,
  28186, 28037, 27524, 26844, 25753, 24219, 22841, 22255, 22180, 22473, 
    22906, 23588, 24591, 25754, 26637, 28029, 27489, 26391, 25801, 25138, 
    24403, 23680,
  28075, 27949, 27395, 26828, 25757, 24311, 22906, 22325, 22139, 22452, 
    22894, 23564, 24717, 25724, 26779, 27862, 27190, 26124, 25671, 25132, 
    24403, 23706,
  27960, 27878, 27339, 26796, 25798, 24359, 22923, 22369, 22168, 22495, 
    22914, 23524, 24460, 25643, 26501, 27764, 27097, 26038, 25554, 25001, 
    24282, 23739,
  27867, 27818, 27293, 26854, 25864, 24448, 22989, 22372, 22200, 22512, 
    22817, 23508, 24445, 25607, 26499, 27650, 27053, 26160, 25671, 25174, 
    24370, 23718,
  27782, 27721, 27217, 26817, 25869, 24538, 23086, 22402, 22208, 22520, 
    22864, 23589, 24504, 25689, 26387, 27529, 27190, 26232, 25747, 25087, 
    24414, 23852,
  27675, 27567, 27020, 26674, 25854, 24574, 23131, 22451, 22240, 22500, 
    22870, 23573, 24536, 25679, 26516, 27097, 26892, 26189, 25732, 25187, 
    24541, 23978,
  27527, 27386, 26723, 26421, 25743, 24540, 23190, 22498, 22251, 22522, 
    22841, 23497, 24447, 25489, 26879, 26429, 25828, 25648, 25450, 25050, 
    24503, 23885,
  27336, 27212, 26548, 26335, 25669, 24644, 23217, 22539, 22245, 22525, 
    22872, 23502, 24402, 25551, 26685, 25919, 24478, 24948, 25050, 24795, 
    24356, 23751,
  27143, 27059, 26563, 26345, 25731, 24646, 23314, 22574, 22286, 22493, 
    22866, 23456, 24242, 25657, 26510, 26220, 25492, 25424, 25264, 24931, 
    24381, 23837,
  27001, 26940, 26712, 26450, 25800, 24727, 23384, 22642, 22347, 22547, 
    22886, 23448, 24342, 25388, 26799, 26609, 26045, 25539, 25270, 24875, 
    24330, 23730,
  26948, 26886, 26743, 26509, 25917, 24766, 23397, 22686, 22355, 22464, 
    22846, 23390, 24310, 25581, 26692, 26687, 25665, 25402, 25153, 24831, 
    24272, 23803,
  26979, 26918, 26778, 26515, 25937, 24836, 23421, 22691, 22355, 22504, 
    22888, 23435, 24377, 25667, 26525, 26846, 26101, 25646, 25332, 24856, 
    24202, 23756,
  27070, 27020, 26867, 26663, 26095, 24934, 23487, 22726, 22369, 22520, 
    22905, 23554, 24428, 25506, 26806, 27123, 26585, 25870, 25462, 24967, 
    24297, 23842,
  27190, 27140, 27047, 26784, 26091, 24951, 23546, 22740, 22384, 22566, 
    22828, 23404, 24504, 25423, 26982, 27310, 26785, 25899, 25386, 24911, 
    24259, 23735,
  27300, 27226, 27075, 26797, 26117, 24970, 23559, 22779, 22366, 22520, 
    22885, 23399, 24152, 25688, 26903, 27304, 26360, 25487, 25151, 24687, 
    24137, 23714,
  27356, 27256, 27069, 26778, 26162, 25018, 23618, 22814, 22427, 22525, 
    22790, 23396, 24314, 25485, 26381, 27218, 26249, 25508, 25193, 24892, 
    24284, 23848,
  27324, 27230, 27035, 26704, 26157, 25049, 23677, 22831, 22465, 22542, 
    22810, 23347, 24328, 25452, 26546, 27246, 26592, 25832, 25365, 24960, 
    24283, 23687,
  27202, 27143, 27010, 26726, 26145, 25088, 23673, 22846, 22459, 22525, 
    22784, 23357, 24348, 25447, 26401, 27249, 26840, 26121, 25632, 25090, 
    24372, 23881,
  27009, 26980, 26985, 26697, 26097, 25057, 23673, 22884, 22500, 22548, 
    22887, 23393, 24217, 25515, 26679, 27257, 26872, 26200, 25681, 25183, 
    24442, 23800,
  26775, 26748, 26985, 26694, 26125, 25079, 23729, 22934, 22491, 22547, 
    22843, 23382, 24254, 25333, 26468, 27154, 26846, 26185, 25729, 25214, 
    24454, 23813,
  26535, 26496, 26745, 26657, 26114, 25149, 23766, 22963, 22552, 22547, 
    22815, 23410, 24347, 25189, 26382, 26990, 26529, 26099, 25681, 25170, 
    24517, 23820,
  26338, 26299, 26765, 26619, 26145, 25151, 23759, 22960, 22537, 22532, 
    22840, 23409, 24281, 25433, 26625, 26960, 26323, 26004, 25673, 25294, 
    24606, 23926,
  26236, 26207, 26724, 26604, 26182, 25160, 23787, 23001, 22580, 22535, 
    22911, 23384, 24334, 25435, 26476, 27107, 26790, 26279, 25866, 25306, 
    24631, 23980,
  26247, 26213, 26762, 26616, 26174, 25148, 23832, 23039, 22560, 22534, 
    22785, 23462, 24164, 25149, 26613, 27228, 27032, 26409, 25963, 25430, 
    24688, 24073,
  26339, 26277, 26835, 26662, 26196, 25120, 23852, 23036, 22589, 22583, 
    22873, 23447, 24219, 25302, 26584, 27204, 26920, 26373, 25997, 25436, 
    24841, 24119,
  26452, 26357, 26790, 26701, 26165, 25190, 23814, 23000, 22551, 22543, 
    22748, 23381, 24253, 25409, 26610, 27119, 26871, 26394, 26051, 25567, 
    24866, 24193,
  26527, 26417, 26754, 26634, 26159, 25199, 23870, 23036, 22621, 22632, 
    22805, 23299, 24127, 25340, 26620, 27110, 26951, 26423, 26004, 25542, 
    24860, 24166,
  26537, 26424, 26787, 26679, 26201, 25271, 23873, 23082, 22641, 22551, 
    22856, 23352, 24280, 25088, 26438, 27170, 27138, 26459, 26059, 25666, 
    24910, 24233,
  26486, 26374, 26792, 26678, 26248, 25237, 23956, 23085, 22576, 22606, 
    22921, 23410, 24185, 25251, 26467, 27242, 27263, 26603, 26072, 25603, 
    24993, 24326,
  26415, 26302, 26739, 26660, 26187, 25263, 23873, 23144, 22623, 22591, 
    22759, 23334, 24225, 25216, 26372, 27178, 27250, 26668, 26217, 25796, 
    25050, 24473,
  26370, 26260, 26675, 26560, 26160, 25201, 23921, 23109, 22655, 22590, 
    22821, 23390, 24020, 25204, 26350, 27089, 27219, 26566, 26210, 25759, 
    25209, 24553,
  26356, 26258, 26619, 26551, 26147, 25229, 23897, 23111, 22669, 22553, 
    22852, 23250, 24183, 25225, 26547, 26997, 27076, 26559, 26182, 25846, 
    25183, 24540,
  26327, 26253, 26663, 26560, 26164, 25212, 23939, 23149, 22678, 22582, 
    22841, 23380, 24239, 25443, 26369, 26975, 27014, 26538, 26134, 25739, 
    25145, 24673,
  26239, 26199, 26571, 26567, 26089, 25231, 23966, 23164, 22722, 22699, 
    22906, 23341, 24180, 25320, 26591, 26857, 26957, 26516, 26085, 25765, 
    25196, 24660,
  26099, 26087, 26507, 26499, 26096, 25229, 23935, 23170, 22698, 22595, 
    22795, 23260, 24096, 25346, 26532, 26744, 26864, 26371, 26092, 25628, 
    25208, 24647,
  25963, 25959, 26454, 26401, 26115, 25198, 23959, 23173, 22751, 22613, 
    22832, 23409, 24101, 25299, 26617, 26568, 26770, 26328, 26037, 25651, 
    25157, 24800,
  25882, 25867, 26241, 26294, 26026, 25195, 23938, 23170, 22724, 22687, 
    22860, 23363, 23953, 25378, 26398, 26401, 26801, 26335, 26057, 25726, 
    25272, 24820,
  25869, 25840, 26348, 26370, 26095, 25195, 23973, 23170, 22745, 22621, 
    22868, 23351, 24201, 25353, 26369, 26390, 26764, 26349, 26016, 25707, 
    25272, 24961,
  25894, 25862, 26431, 26394, 26110, 25203, 23952, 23202, 22754, 22661, 
    22909, 23371, 24167, 25129, 26495, 26390, 26676, 26270, 25926, 25626, 
    25227, 24894,
  25914, 25898, 26382, 26385, 26081, 25250, 23993, 23252, 22745, 22641, 
    22945, 23313, 24201, 25278, 26710, 26340, 26676, 26248, 25960, 25646, 
    25131, 24807,
  25931, 25937, 26340, 26394, 26089, 25265, 23996, 23234, 22771, 22641, 
    22914, 23313, 24174, 25389, 26226, 26226, 26820, 26349, 25913, 25577, 
    25157, 24806,
  25994, 26014, 26326, 26394, 26141, 25262, 23983, 23196, 22774, 22698, 
    22882, 23355, 24157, 25399, 26810, 26106, 26807, 26298, 25899, 25422, 
    25010, 24652,
  26126, 26151, 26482, 26513, 26209, 25270, 23976, 23213, 22768, 22580, 
    22837, 23376, 24260, 25329, 26604, 26229, 26770, 26234, 25781, 25422, 
    24953, 24505,
  26264, 26290, 26785, 26734, 26272, 25256, 24000, 23199, 22768, 22644, 
    22845, 23350, 24303, 25315, 26121, 26672, 26839, 26241, 25781, 25390, 
    24831, 24552,
  26304, 26333, 26896, 26809, 26292, 25329, 24004, 23199, 22806, 22687, 
    22977, 23386, 24167, 25103, 26337, 26900, 27050, 26254, 25754, 25285, 
    24774, 24398,
  26205, 26242, 26776, 26693, 26284, 25295, 24024, 23207, 22815, 22681, 
    22860, 23241, 24021, 25436, 26490, 26847, 27013, 26320, 25774, 25353, 
    24793, 24418,
  26026, 26082, 26523, 26499, 26181, 25262, 23989, 23246, 22818, 22684, 
    22817, 23363, 24332, 25177, 26349, 26524, 26839, 26313, 25740, 25247, 
    24736, 24418,
  25884, 25960, 26365, 26413, 26092, 25279, 23972, 23207, 22821, 22747, 
    22874, 23317, 24065, 25368, 26622, 26265, 26496, 25995, 25567, 25166, 
    24621, 24190,
  25866, 25944, 26479, 26462, 26154, 25253, 24011, 23240, 22806, 22652, 
    22982, 23345, 24021, 25366, 26457, 26401, 26415, 25865, 25436, 25110, 
    24641, 24244,
  25973, 26035, 26657, 26560, 26184, 25281, 23986, 23269, 22791, 22692, 
    22857, 23279, 24236, 25243, 26685, 26626, 26651, 26075, 25588, 25260, 
    24628, 24257,
  26121, 26177, 26785, 26618, 26221, 25290, 23952, 23222, 22824, 22687, 
    22894, 23318, 24325, 25177, 26687, 26831, 27019, 26363, 25919, 25384, 
    24749, 24277,
  26197, 26279, 26731, 26604, 26224, 25279, 23972, 23222, 22815, 22666, 
    22905, 23460, 24085, 25348, 26235, 26832, 27181, 26660, 26132, 25552, 
    24730, 24231,
  26123, 26250, 26644, 26504, 26141, 25268, 23993, 23252, 22833, 22715, 
    22900, 23350, 24196, 25387, 26809, 26716, 27150, 26696, 26168, 25559, 
    24761, 24264,
  25864, 26017, 26504, 26504, 26129, 25234, 23976, 23219, 22824, 22733, 
    22911, 23340, 24086, 25150, 26575, 26591, 27206, 26760, 26182, 25607, 
    24851, 24257,
  25396, 25540, 26396, 26443, 26138, 25212, 23983, 23222, 22786, 22744, 
    22900, 23325, 24379, 25264, 26782, 26476, 27113, 26754, 26209, 25632, 
    24876, 24298,
  24686, 24812, 26056, 26235, 26041, 25155, 23948, 23217, 22871, 22764, 
    22997, 23353, 24204, 25420, 26425, 26134, 27013, 26804, 26251, 25770, 
    24947, 24324,
  23721, 23866, 25561, 25917, 25918, 25139, 23945, 23173, 22824, 22730, 
    22960, 23331, 24105, 25389, 26435, 25493, 26770, 26819, 26389, 25776, 
    25099, 24492,
  22560, 22775, 25039, 25578, 25734, 25116, 23900, 23217, 22830, 22721, 
    22946, 23311, 24266, 25402, 26579, 24880, 26528, 26862, 26417, 25851, 
    25093, 24485,
  21362, 21670, 24456, 25220, 25560, 25052, 23917, 23229, 22827, 22788, 
    22906, 23387, 24054, 25292, 26270, 24393, 26428, 26740, 26313, 25764, 
    25062, 24439,
  20361, 20738, 23586, 24606, 25322, 24951, 23903, 23235, 22842, 22719, 
    23023, 23476, 24113, 25227, 26384, 23370, 25649, 26559, 26334, 25726, 
    25049, 24412,
  19790, 20184, 22967, 24237, 25131, 24900, 23924, 23182, 22851, 22779, 
    22952, 23382, 24276, 25294, 26407, 22560, 25176, 26588, 26334, 25864, 
    25100, 24459,
  19762, 20127, 23282, 24393, 25173, 24929, 23851, 23214, 22816, 22831, 
    23000, 23400, 24155, 25239, 26469, 22883, 25593, 26566, 26341, 25826, 
    25120, 24593,
  20197, 20500, 23845, 24711, 25268, 24895, 23869, 23217, 22892, 22782, 
    22964, 23463, 24230, 25309, 26488, 23478, 25787, 26603, 26376, 25901, 
    25177, 24607,
  20851, 21073, 24167, 24924, 25354, 24878, 23841, 23218, 22887, 22840, 
    22938, 23408, 24351, 25360, 26513, 23868, 25781, 26617, 26376, 25870, 
    25145, 24714,
  21450, 21608, 24332, 25110, 25414, 24915, 23841, 23232, 22860, 22817, 
    22987, 23385, 24292, 25488, 26719, 24177, 25968, 26654, 26307, 25896, 
    25222, 24647,
  21842, 21981, 24350, 25054, 25369, 24859, 23814, 23189, 22933, 22840, 
    23075, 23421, 24309, 25332, 26321, 24182, 25893, 26646, 26314, 25826, 
    25222, 24708,
  22035, 22187, 24297, 25016, 25374, 24910, 23814, 23177, 22884, 22869, 
    23004, 23469, 24154, 25265, 26700, 24098, 25825, 26567, 26231, 25840, 
    25139, 24607,
  22108, 22257, 24292, 24984, 25357, 24851, 23828, 23168, 22872, 22838, 
    22993, 23423, 24181, 25396, 26674, 23975, 25706, 26538, 26259, 25747, 
    25082, 24574,
  22111, 22217, 24376, 25005, 25338, 24800, 23779, 23192, 22864, 22890, 
    23067, 23538, 24346, 25396, 26529, 24067, 25676, 26445, 26121, 25710, 
    25063, 24594,
  22031, 22096, 24520, 25127, 25355, 24814, 23779, 23186, 22885, 22867, 
    23056, 23436, 24418, 25570, 27010, 24387, 26049, 26531, 26232, 25679, 
    25064, 24688,
  21861, 21940, 24545, 25138, 25346, 24809, 23724, 23163, 22855, 22853, 
    23094, 23460, 24300, 25363, 26707, 24601, 26168, 26501, 26218, 25629, 
    25140, 24649,
  21653, 21799, 24249, 25014, 25264, 24700, 23703, 23139, 22859, 22839, 
    23122, 23439, 24350, 25678, 26496, 24384, 26054, 26553, 26149, 25835, 
    25134, 24669,
  21490, 21701, 24004, 24874, 25238, 24717, 23686, 23146, 22885, 22819, 
    23060, 23572, 24391, 25405, 26972, 24091, 25962, 26429, 26129, 25785, 
    25160, 24656,
  21397, 21640, 24125, 24912, 25221, 24728, 23718, 23143, 22889, 22868, 
    23006, 23516, 24315, 25471, 26497, 24118, 25987, 26401, 26135, 25754, 
    25147, 24649,
  21300, 21565, 24348, 25052, 25261, 24647, 23680, 23131, 22851, 22862, 
    23117, 23481, 24370, 25584, 26629, 24394, 26074, 26373, 25984, 25642, 
    25084, 24522,
  21080, 21383, 24460, 25103, 25273, 24647, 23645, 23117, 22895, 22889, 
    23163, 23545, 24515, 25606, 26860, 24449, 26062, 26374, 26060, 25660, 
    24989, 24603,
  20675, 21020, 24123, 24929, 25249, 24661, 23635, 23103, 22895, 22883, 
    23041, 23512, 24378, 25615, 26667, 24100, 25994, 26410, 26047, 25649, 
    25072, 24637,
  20164, 20510, 23753, 24756, 25161, 24569, 23611, 23085, 22927, 22866, 
    23030, 23507, 24395, 25722, 26866, 23520, 25869, 26359, 25999, 25631, 
    25078, 24590,
  19754, 20034, 23553, 24646, 25087, 24547, 23576, 23076, 22896, 22946, 
    23124, 23599, 24368, 25371, 26509, 23099, 25657, 26324, 25972, 25531, 
    25015, 24463,
  19666, 19833, 23665, 24700, 25059, 24516, 23521, 23130, 22896, 22932, 
    23061, 23523, 24366, 25732, 26728, 22968, 25609, 26287, 25929, 25519, 
    24952, 24323,
  20008, 20056, 23675, 24692, 25130, 24511, 23532, 23091, 22948, 22899, 
    23155, 23558, 24595, 25888, 26851, 22919, 25497, 26207, 25924, 25557, 
    24964, 24350,
  20701, 20667, 23974, 24811, 25039, 24418, 23556, 23048, 22902, 22924, 
    23122, 23576, 24490, 25706, 26829, 23117, 25634, 26301, 26006, 25632, 
    25105, 24438,
  21533, 21473, 24466, 25045, 25136, 24438, 23490, 23033, 22847, 22905, 
    23162, 23597, 24620, 25726, 26867, 23814, 25882, 26360, 26076, 25762, 
    25131, 24625,
  22275, 22229, 24834, 25193, 25131, 24377, 23442, 23034, 22935, 22902, 
    23091, 23666, 24520, 25767, 26829, 24368, 26095, 26267, 26021, 25676, 
    25144, 24759,
  22788, 22765, 24923, 25296, 25168, 24369, 23394, 23057, 22915, 23003, 
    23100, 23633, 24448, 26021, 27032, 24524, 25970, 26216, 25951, 25663, 
    25029, 24605,
  23077, 23067, 24992, 25312, 25091, 24318, 23422, 23058, 22971, 22986, 
    23023, 23684, 24528, 25816, 26857, 24446, 26088, 26238, 25959, 25645, 
    25042, 24586,
  23241, 23240, 25078, 25339, 25091, 24299, 23366, 23046, 22933, 22975, 
    23180, 23687, 24518, 25751, 26810, 24420, 26064, 26239, 25882, 25732, 
    25005, 24506,
  23386, 23383, 25134, 25337, 25042, 24204, 23384, 23017, 22939, 22989, 
    23214, 23649, 24533, 25860, 27003, 24467, 26064, 26224, 25891, 25601, 
    24967, 24399,
  23573, 23535, 25207, 25353, 25049, 24201, 23360, 23008, 22968, 23033, 
    23226, 23748, 24649, 26085, 26816, 24547, 26057, 26109, 25822, 25534, 
    24878, 24399,
  23817, 23725, 25347, 25396, 24963, 24128, 23319, 23041, 22939, 22976, 
    23167, 23776, 24610, 25898, 27013, 24550, 26107, 26124, 25835, 25404, 
    24796, 24213,
  24072, 23952, 25395, 25412, 24951, 24067, 23316, 23050, 22948, 22950, 
    23201, 23754, 24785, 26001, 27154, 24625, 26046, 26103, 25754, 25373, 
    24847, 24220,
  24198, 24088, 25403, 25423, 24883, 24051, 23257, 22994, 22963, 23045, 
    23164, 23706, 24840, 26059, 27260, 24658, 26065, 25966, 25629, 25311, 
    24701, 24167,
  24065, 23956, 25461, 25388, 24829, 23911, 23247, 22992, 23001, 23025, 
    23273, 23838, 24704, 26029, 26954, 24789, 26051, 25894, 25499, 25094, 
    24536, 24093,
  23767, 23625, 25489, 25362, 24778, 23883, 23184, 22995, 22961, 23054, 
    23279, 23803, 24771, 26026, 27290, 24797, 26096, 25815, 25410, 25020, 
    24390, 24074,
  23610, 23443, 25492, 25316, 24686, 23816, 23153, 22998, 22970, 23026, 
    23194, 23816, 24917, 26245, 27009, 24707, 26090, 25714, 25397, 24984, 
    24365, 23954,
  28133, 28000, 27450, 26838, 25596, 24094, 22735, 22231, 22151, 22487, 
    22805, 23637, 24804, 25841, 26429, 28032, 27354, 26445, 25894, 25280, 
    24406, 23703,
  28078, 27946, 27364, 26792, 25668, 24180, 22773, 22287, 22139, 22446, 
    22873, 23475, 24580, 25562, 26537, 27792, 26931, 26192, 25728, 25174, 
    24362, 23763,
  27956, 27836, 27254, 26709, 25691, 24351, 22891, 22340, 22142, 22440, 
    22819, 23574, 24637, 25574, 26563, 27543, 26726, 25969, 25542, 25037, 
    24406, 23730,
  27837, 27751, 27154, 26654, 25765, 24427, 22981, 22331, 22192, 22480, 
    22926, 23531, 24530, 25511, 26815, 27443, 26787, 25925, 25452, 24975, 
    24374, 23716,
  27749, 27701, 27169, 26714, 25819, 24466, 23033, 22434, 22259, 22500, 
    22929, 23518, 24498, 25820, 26670, 27387, 26800, 26032, 25624, 25136, 
    24456, 23796,
  27678, 27631, 27070, 26660, 25832, 24538, 23095, 22460, 22217, 22485, 
    22909, 23520, 24569, 25666, 26747, 27214, 26906, 26141, 25693, 25148, 
    24481, 23862,
  27604, 27511, 26819, 26493, 25767, 24569, 23146, 22462, 22234, 22479, 
    22897, 23593, 24510, 25618, 26560, 26723, 26364, 25924, 25555, 25036, 
    24424, 23848,
  27510, 27366, 26700, 26375, 25713, 24549, 23237, 22498, 22266, 22479, 
    22882, 23364, 24463, 25631, 26557, 26198, 24984, 25175, 25093, 24844, 
    24340, 23848,
  27382, 27231, 26664, 26420, 25775, 24624, 23264, 22551, 22254, 22490, 
    22856, 23453, 24315, 25503, 26409, 26215, 24635, 24836, 24879, 24700, 
    24251, 23794,
  27227, 27114, 26775, 26479, 25847, 24677, 23313, 22580, 22327, 22467, 
    22845, 23346, 24346, 25480, 26747, 26642, 26078, 25592, 25354, 24898, 
    24327, 23860,
  27083, 27010, 26829, 26503, 25864, 24776, 23354, 22650, 22321, 22478, 
    22816, 23463, 24405, 25431, 26523, 26860, 26438, 25779, 25437, 24923, 
    24333, 23867,
  26990, 26936, 26851, 26535, 25938, 24753, 23440, 22664, 22364, 22526, 
    22784, 23404, 24307, 25591, 26507, 26897, 26246, 25794, 25423, 24911, 
    24390, 23840,
  26968, 26920, 26869, 26554, 25926, 24845, 23468, 22732, 22376, 22540, 
    22878, 23472, 24361, 25456, 26671, 26953, 26401, 25887, 25485, 24972, 
    24364, 23846,
  27019, 26973, 26912, 26604, 26026, 24926, 23482, 22750, 22332, 22531, 
    22847, 23439, 24328, 25751, 26528, 27139, 26818, 26139, 25629, 25003, 
    24377, 23793,
  27122, 27067, 26973, 26737, 26078, 24926, 23520, 22755, 22399, 22477, 
    22832, 23446, 24390, 25414, 26564, 27257, 26867, 26016, 25491, 24990, 
    24344, 23839,
  27232, 27153, 27079, 26775, 26115, 25030, 23571, 22820, 22413, 22596, 
    22821, 23410, 24195, 25567, 26887, 27279, 26556, 25785, 25422, 24897, 
    24319, 23805,
  27295, 27196, 27001, 26791, 26160, 25018, 23651, 22834, 22448, 22548, 
    22903, 23504, 24298, 25532, 26542, 27263, 26556, 25959, 25546, 25002, 
    24287, 23812,
  27270, 27180, 27007, 26737, 26140, 24990, 23623, 22872, 22459, 22481, 
    22766, 23346, 24206, 25348, 26598, 27244, 26842, 26260, 25759, 25226, 
    24483, 23878,
  27147, 27092, 26988, 26720, 26129, 25063, 23716, 22887, 22532, 22570, 
    22794, 23448, 24286, 25506, 26794, 27146, 26854, 26282, 25779, 25325, 
    24515, 23878,
  26943, 26911, 26879, 26675, 26085, 25021, 23702, 22942, 22497, 22538, 
    22805, 23414, 24243, 25448, 26406, 27024, 26549, 26151, 25807, 25349, 
    24553, 24085,
  26693, 26652, 26803, 26589, 26054, 25090, 23723, 22933, 22514, 22506, 
    22828, 23397, 24270, 25497, 26384, 26965, 26444, 26123, 25834, 25349, 
    24667, 24038,
  26440, 26381, 26724, 26570, 26091, 25068, 23699, 22936, 22508, 22538, 
    22887, 23404, 24312, 25294, 26670, 26965, 26456, 26151, 25799, 25361, 
    24762, 24098,
  26240, 26182, 26632, 26543, 26106, 25130, 23761, 22977, 22519, 22543, 
    22899, 23480, 24321, 25217, 26401, 27041, 26854, 26347, 25951, 25498, 
    24781, 24178,
  26136, 26098, 26732, 26589, 26134, 25152, 23768, 22997, 22543, 22494, 
    22827, 23350, 24193, 25464, 26692, 27099, 26978, 26498, 26041, 25647, 
    24902, 24278,
  26132, 26102, 26716, 26623, 26179, 25166, 23809, 22977, 22549, 22540, 
    22918, 23378, 24249, 25280, 26493, 27116, 27047, 26491, 26068, 25560, 
    24882, 24218,
  26189, 26135, 26632, 26612, 26160, 25168, 23792, 23056, 22577, 22554, 
    22841, 23299, 24163, 25347, 26599, 27122, 27065, 26520, 26101, 25628, 
    24965, 24371,
  26251, 26155, 26635, 26521, 26171, 25182, 23854, 23047, 22630, 22525, 
    22852, 23337, 24066, 25247, 26524, 27019, 27059, 26576, 26232, 25765, 
    25079, 24378,
  26282, 26153, 26541, 26545, 26188, 25162, 23878, 23056, 22641, 22590, 
    22880, 23362, 24175, 25161, 26747, 26924, 27003, 26534, 26164, 25657, 
    25009, 24404,
  26272, 26133, 26531, 26515, 26166, 25241, 23889, 23076, 22670, 22567, 
    22920, 23341, 24103, 25263, 26150, 26926, 27207, 26591, 26178, 25671, 
    25028, 24424,
  26240, 26109, 26526, 26582, 26214, 25210, 23906, 23061, 22694, 22619, 
    22834, 23407, 24222, 25217, 26635, 26939, 27251, 26562, 26226, 25807, 
    25225, 24585,
  26228, 26115, 26560, 26579, 26174, 25241, 23937, 23070, 22661, 22627, 
    22854, 23422, 24217, 25282, 26497, 26960, 27226, 26728, 26309, 25907, 
    25212, 24591,
  26280, 26190, 26528, 26531, 26139, 25213, 23919, 23105, 22696, 22636, 
    22842, 23374, 24165, 25119, 26609, 26926, 27132, 26620, 26309, 25882, 
    25231, 24779,
  26395, 26337, 26607, 26612, 26128, 25176, 23902, 23152, 22688, 22653, 
    22899, 23267, 24167, 25065, 26570, 26925, 26922, 26554, 26212, 25857, 
    25288, 24805,
  26519, 26500, 26792, 26617, 26135, 25218, 23922, 23137, 22640, 22635, 
    22862, 23310, 24233, 25261, 26441, 26979, 26828, 26475, 26176, 25820, 
    25320, 24772,
  26588, 26605, 26756, 26631, 26113, 25184, 23915, 23140, 22725, 22621, 
    22796, 23282, 24253, 25261, 26621, 26945, 26828, 26439, 26107, 25713, 
    25276, 24932,
  26579, 26618, 26870, 26644, 26176, 25212, 23937, 23119, 22719, 22638, 
    22859, 23325, 24031, 25258, 26198, 26919, 26810, 26388, 25976, 25720, 
    25275, 24791,
  26523, 26572, 26764, 26671, 26142, 25243, 23954, 23190, 22716, 22638, 
    22842, 23325, 24208, 25274, 26453, 26851, 26878, 26257, 25915, 25651, 
    25263, 24892,
  26474, 26524, 26748, 26635, 26153, 25229, 23964, 23187, 22783, 22621, 
    22881, 23383, 24136, 25265, 26489, 26766, 26840, 26338, 25949, 25719, 
    25294, 24925,
  26467, 26513, 26799, 26695, 26176, 25226, 23957, 23207, 22713, 22615, 
    22793, 23403, 24245, 25360, 26499, 26807, 26803, 26316, 25982, 25663, 
    25211, 24919,
  26495, 26535, 26870, 26635, 26185, 25192, 23988, 23210, 22748, 22609, 
    22836, 23393, 24164, 25276, 26535, 26831, 26728, 26200, 25866, 25545, 
    25084, 24818,
  26524, 26562, 26776, 26700, 26210, 25248, 23967, 23190, 22745, 22615, 
    23004, 23367, 24045, 25272, 26475, 26800, 26790, 26193, 25797, 25508, 
    25058, 24697,
  26539, 26578, 26797, 26728, 26190, 25231, 23971, 23184, 22768, 22632, 
    22867, 23421, 24178, 25418, 26432, 26679, 26822, 26099, 25707, 25327, 
    24912, 24529,
  26555, 26595, 26792, 26679, 26229, 25254, 24033, 23222, 22763, 22651, 
    22841, 23431, 24218, 25388, 26421, 26629, 26210, 25593, 25313, 25084, 
    24663, 24449,
  26569, 26611, 26982, 26784, 26239, 25296, 23988, 23222, 22812, 22680, 
    22855, 23360, 24292, 25451, 26798, 26719, 25657, 25081, 24968, 24767, 
    24459, 24274,
  26520, 26570, 26882, 26859, 26229, 25307, 23970, 23222, 22800, 22646, 
    22861, 23388, 24225, 25411, 26579, 26842, 26068, 25442, 25155, 24904, 
    24548, 24161,
  26348, 26408, 26814, 26684, 26248, 25271, 24005, 23246, 22786, 22686, 
    22878, 23301, 24097, 25479, 26554, 26800, 26235, 25607, 25306, 24966, 
    24516, 24207,
  26074, 26138, 26464, 26509, 26116, 25228, 23977, 23219, 22771, 22703, 
    22938, 23393, 24257, 25388, 26373, 26514, 26460, 25947, 25520, 25072, 
    24599, 24355,
  25808, 25869, 26354, 26379, 26132, 25254, 23960, 23207, 22783, 22729, 
    23020, 23390, 24171, 25479, 26639, 26271, 26398, 25932, 25479, 25134, 
    24593, 24187,
  25667, 25724, 26228, 26323, 26087, 25226, 23998, 23243, 22789, 22712, 
    22972, 23395, 24158, 25309, 26582, 26040, 26310, 25982, 25486, 25078, 
    24612, 24187,
  25708, 25761, 26238, 26350, 26087, 25251, 23974, 23240, 22836, 22740, 
    23015, 23398, 24227, 25045, 26819, 26185, 26547, 26171, 25721, 25165, 
    24708, 24207,
  25893, 25943, 26509, 26568, 26213, 25265, 23998, 23252, 22800, 22706, 
    22909, 23365, 24299, 25534, 27057, 26551, 26915, 26395, 25976, 25383, 
    24784, 24254,
  26111, 26166, 26768, 26706, 26248, 25251, 23974, 23213, 22830, 22732, 
    22910, 23360, 24220, 25516, 26426, 26875, 27257, 26640, 26121, 25563, 
    24873, 24442,
  26239, 26309, 26819, 26719, 26248, 25282, 24012, 23237, 22836, 22740, 
    22904, 23367, 24207, 25481, 26567, 26937, 27382, 26749, 26218, 25607, 
    24956, 24489,
  26192, 26281, 26649, 26671, 26225, 25282, 23984, 23210, 22818, 22764, 
    22995, 23469, 24333, 25430, 26788, 26806, 27345, 26800, 26239, 25737, 
    24950, 24442,
  25927, 26032, 26520, 26550, 26132, 25276, 23967, 23243, 22839, 22740, 
    22952, 23433, 24237, 25388, 26579, 26601, 27121, 26771, 26246, 25806, 
    25039, 24623,
  25410, 25530, 26391, 26445, 26132, 25212, 23953, 23240, 22830, 22740, 
    23058, 23454, 24255, 25374, 26491, 26485, 27164, 26843, 26363, 25757, 
    25103, 24529,
  24616, 24763, 26260, 26364, 26067, 25240, 23985, 23225, 22898, 22767, 
    22967, 23347, 24272, 25460, 26363, 26279, 27171, 26885, 26418, 25769, 
    25115, 24664,
  23570, 23771, 25764, 26025, 25953, 25164, 23929, 23178, 22812, 22784, 
    22910, 23413, 24368, 25320, 26912, 25757, 26996, 26879, 26376, 25906, 
    25185, 24583,
  22388, 22667, 24935, 25515, 25666, 25097, 23954, 23213, 22848, 22784, 
    23024, 23419, 24048, 25346, 26501, 24961, 26498, 26713, 26329, 25794, 
    25141, 24550,
  21272, 21622, 24166, 24968, 25467, 25016, 23905, 23175, 22874, 22770, 
    23007, 23470, 24356, 25372, 26414, 24007, 26031, 26604, 26301, 25862, 
    25193, 24550,
  20451, 20829, 23355, 24527, 25198, 24957, 23895, 23243, 22842, 22830, 
    22982, 23365, 24236, 25333, 26729, 23062, 25383, 26612, 26384, 25826, 
    25078, 24490,
  20090, 20450, 23157, 24338, 25172, 24943, 23888, 23241, 22848, 22870, 
    23013, 23437, 24359, 25370, 26210, 22670, 25240, 26510, 26349, 25838, 
    25250, 24610,
  20223, 20537, 23477, 24532, 25255, 24937, 23864, 23226, 22874, 22848, 
    22999, 23480, 24201, 25263, 27017, 23134, 25520, 26612, 26398, 25981, 
    25218, 24658,
  20719, 20969, 23994, 24789, 25347, 24890, 23843, 23176, 22910, 22807, 
    22996, 23561, 24268, 25191, 26521, 23727, 25776, 26612, 26370, 25913, 
    25295, 24638,
  21333, 21509, 24355, 25041, 25372, 24938, 23916, 23205, 22843, 22879, 
    23045, 23526, 24268, 25454, 26864, 24189, 26000, 26641, 26385, 25913, 
    25301, 24725,
  21830, 21951, 24390, 25058, 25389, 24882, 23829, 23229, 22843, 22848, 
    23116, 23481, 24357, 25691, 26844, 24225, 25925, 26591, 26392, 25957, 
    25346, 24873,
  22108, 22217, 24316, 25012, 25364, 24898, 23857, 23203, 22875, 22886, 
    23022, 23503, 24377, 25660, 26609, 24021, 25645, 26598, 26343, 25889, 
    25206, 24712,
  22205, 22324, 24355, 24988, 25370, 24857, 23795, 23174, 22846, 22929, 
    23062, 23552, 24207, 25300, 26499, 24043, 25720, 26519, 26198, 25746, 
    25181, 24739,
  22200, 22307, 24334, 25012, 25347, 24874, 23784, 23192, 22922, 22877, 
    23091, 23562, 24325, 25570, 26691, 24010, 25720, 26519, 26212, 25746, 
    25130, 24672,
  22118, 22185, 24418, 25056, 25333, 24773, 23774, 23153, 22876, 22898, 
    23023, 23454, 24311, 25456, 26754, 24179, 25895, 26476, 26164, 25751, 
    25092, 24646,
  21932, 21980, 24497, 25115, 25353, 24762, 23785, 23166, 22908, 22892, 
    23140, 23436, 24311, 25489, 26616, 24502, 26119, 26504, 26185, 25721, 
    25124, 24659,
  21652, 21736, 24200, 24937, 25236, 24720, 23698, 23139, 22870, 22910, 
    23089, 23423, 24392, 25464, 26929, 24385, 26038, 26491, 26137, 25684, 
    25169, 24746,
  21370, 21524, 23886, 24760, 25204, 24694, 23678, 23142, 22844, 22896, 
    23101, 23545, 24378, 25559, 26687, 23961, 25832, 26498, 26137, 25728, 
    25137, 24814,
  21214, 21415, 23735, 24682, 25170, 24701, 23685, 23125, 22868, 22878, 
    23101, 23528, 24376, 25654, 26732, 23821, 25739, 26419, 26144, 25740, 
    25214, 24734,
  21232, 21442, 23945, 24752, 25179, 24675, 23685, 23128, 22895, 22919, 
    23104, 23622, 24346, 25515, 26612, 23974, 25807, 26404, 26082, 25728, 
    25221, 24754,
  21337, 21559, 24308, 25005, 25268, 24637, 23699, 23099, 22889, 22939, 
    23081, 23516, 24462, 25483, 26643, 24381, 26057, 26360, 26097, 25641, 
    25170, 24794,
  21369, 21643, 24465, 25078, 25274, 24600, 23647, 23096, 22874, 22916, 
    23093, 23658, 24440, 25695, 26760, 24612, 26238, 26419, 26062, 25754, 
    25221, 24641,
  21226, 21566, 24450, 25043, 25208, 24645, 23619, 23137, 22922, 22986, 
    23147, 23666, 24236, 25674, 26806, 24477, 26164, 26412, 26042, 25648, 
    25151, 24681,
  20946, 21305, 24146, 24955, 25202, 24598, 23599, 23126, 22896, 22948, 
    23185, 23608, 24485, 25546, 26879, 24026, 25965, 26369, 26056, 25642, 
    25152, 24601,
  20686, 20987, 24093, 24909, 25157, 24539, 23610, 23097, 22887, 23014, 
    23065, 23697, 24397, 25756, 26950, 23763, 25685, 26304, 25951, 25635, 
    25025, 24414,
  20622, 20812, 24179, 24941, 25131, 24522, 23568, 23103, 22911, 23006, 
    23120, 23652, 24530, 25623, 26585, 23729, 25853, 26326, 25966, 25654, 
    24987, 24461,
  20841, 20917, 24281, 24952, 25148, 24450, 23537, 23079, 22934, 22992, 
    23214, 23659, 24506, 25676, 26932, 23651, 25791, 26341, 26056, 25693, 
    25082, 24562,
  21299, 21298, 24357, 25044, 25177, 24475, 23517, 23068, 22897, 23012, 
    23114, 23756, 24570, 25870, 27054, 23709, 25822, 26334, 26043, 25687, 
    25178, 24609,
  21862, 21836, 24623, 25138, 25146, 24464, 23482, 23115, 22955, 23025, 
    23274, 23536, 24607, 26004, 26685, 24060, 25996, 26298, 26091, 25804, 
    25172, 24689,
  22383, 22372, 24854, 25246, 25152, 24422, 23475, 23083, 22909, 22999, 
    23155, 23614, 24595, 25857, 26965, 24355, 26040, 26313, 26057, 25718, 
    25236, 24690,
  22772, 22788, 24908, 25287, 25169, 24341, 23440, 23080, 22956, 22985, 
    23220, 23668, 24546, 25742, 27129, 24396, 25860, 26334, 26071, 25718, 
    25128, 24670,
  23030, 23065, 24984, 25276, 25069, 24316, 23430, 23063, 22947, 23062, 
    23118, 23668, 24775, 26094, 26674, 24399, 25960, 26291, 26009, 25694, 
    25090, 24630,
  23221, 23263, 25012, 25360, 25043, 24280, 23393, 23072, 22968, 22983, 
    23176, 23610, 24470, 25831, 27125, 24435, 26015, 26234, 25913, 25563, 
    25072, 24577,
  23409, 23438, 25134, 25395, 25061, 24219, 23376, 23081, 22963, 23043, 
    23161, 23704, 24692, 25996, 27215, 24481, 26035, 26321, 25968, 25526, 
    25002, 24410,
  23632, 23615, 25212, 25357, 24981, 24236, 23358, 23067, 22948, 23029, 
    23188, 23689, 24769, 25947, 27010, 24531, 26066, 26154, 25851, 25545, 
    25002, 24491,
  23903, 23822, 25308, 25395, 24949, 24115, 23310, 23017, 22989, 23044, 
    23225, 23786, 24677, 25943, 27106, 24573, 26147, 26154, 25885, 25446, 
    24926, 24451,
  24182, 24060, 25403, 25425, 24907, 24076, 23269, 23038, 22948, 23107, 
    23216, 23802, 24747, 26079, 27326, 24609, 26022, 26069, 25810, 25304, 
    24838, 24337,
  24325, 24208, 25403, 25382, 24907, 24015, 23289, 23047, 23016, 23012, 
    23197, 23743, 24851, 25990, 27167, 24698, 26016, 26082, 25749, 25285, 
    24787, 24304,
  24202, 24099, 25481, 25382, 24876, 23940, 23255, 23009, 22978, 23001, 
    23265, 23797, 24821, 26062, 27310, 24828, 25967, 25868, 25577, 25187, 
    24615, 24137,
  23908, 23795, 25446, 25353, 24810, 23900, 23207, 23056, 23026, 23030, 
    23266, 23835, 24725, 26054, 26772, 24884, 26110, 25868, 25487, 25007, 
    24495, 24057,
  23751, 23627, 25436, 25280, 24705, 23850, 23179, 22998, 22952, 23022, 
    23192, 23970, 24829, 26218, 27293, 24772, 26110, 25767, 25377, 24908, 
    24457, 23971,
  28044, 27942, 27354, 26734, 25594, 24116, 22755, 22263, 22132, 22492, 
    22878, 23636, 24497, 25749, 26472, 27882, 27268, 26260, 25726, 25136, 
    24258, 23554,
  27988, 27884, 27234, 26663, 25694, 24183, 22824, 22266, 22149, 22555, 
    22904, 23605, 24740, 25835, 27060, 27573, 26907, 26044, 25582, 25011, 
    24347, 23734,
  27865, 27765, 27165, 26554, 25634, 24266, 22911, 22354, 22135, 22589, 
    22940, 23650, 24642, 25646, 26797, 27322, 26645, 25965, 25526, 25030, 
    24410, 23881,
  27751, 27677, 27016, 26553, 25676, 24392, 22969, 22365, 22196, 22557, 
    22889, 23589, 24326, 25937, 26682, 27219, 26695, 26022, 25616, 25085, 
    24436, 24001,
  27673, 27636, 26976, 26539, 25703, 24429, 23021, 22430, 22207, 22511, 
    22934, 23548, 24658, 25547, 27095, 27012, 26732, 26094, 25663, 25234, 
    24479, 23927,
  27617, 27587, 26857, 26496, 25722, 24507, 23101, 22453, 22230, 22533, 
    22883, 23571, 24500, 25539, 26763, 26735, 26203, 25748, 25477, 25079, 
    24435, 23867,
  27572, 27497, 26751, 26428, 25728, 24526, 23138, 22497, 22241, 22496, 
    22905, 23543, 24611, 25765, 27116, 26418, 25575, 25539, 25277, 24992, 
    24390, 23900,
  27520, 27388, 26789, 26445, 25782, 24613, 23187, 22517, 22297, 22501, 
    22842, 23507, 24473, 25523, 26847, 26356, 24803, 25041, 25070, 24799, 
    24326, 23866,
  27439, 27290, 26840, 26544, 25799, 24658, 23273, 22538, 22270, 22495, 
    22862, 23550, 24487, 25657, 26560, 26635, 25649, 25423, 25180, 24823, 
    24364, 23866,
  27315, 27200, 26926, 26609, 25873, 24663, 23305, 22606, 22264, 22492, 
    22879, 23539, 24509, 25474, 26862, 26999, 26482, 25840, 25380, 24947, 
    24261, 23845,
  27173, 27106, 26926, 26614, 25928, 24688, 23377, 22623, 22346, 22598, 
    22884, 23425, 24374, 25613, 26241, 27125, 26526, 25747, 25324, 24854, 
    24230, 23872,
  27050, 27018, 26934, 26619, 25932, 24805, 23422, 22667, 22351, 22569, 
    22898, 23519, 24469, 25557, 26731, 27125, 26507, 25804, 25414, 24922, 
    24394, 23878,
  26983, 26965, 26882, 26632, 25954, 24839, 23435, 22746, 22401, 22583, 
    22790, 23493, 24383, 25524, 26663, 27139, 26700, 25940, 25503, 24971, 
    24324, 23871,
  26992, 26972, 26890, 26648, 26022, 24926, 23515, 22749, 22394, 22502, 
    22915, 23396, 24259, 25594, 26507, 27206, 27042, 26200, 25682, 25145, 
    24457, 24018,
  27068, 27029, 26918, 26713, 26032, 24951, 23522, 22766, 22409, 22533, 
    22812, 23365, 24404, 25640, 26825, 27285, 27079, 26357, 25765, 25213, 
    24476, 23897,
  27168, 27100, 26960, 26713, 26025, 24945, 23563, 22810, 22449, 22593, 
    22849, 23418, 24242, 25607, 26647, 27293, 27079, 26401, 25889, 25231, 
    24463, 23810,
  27229, 27151, 27051, 26745, 26129, 24970, 23629, 22863, 22508, 22573, 
    22957, 23497, 24382, 25442, 26468, 27234, 27092, 26373, 25901, 25274, 
    24501, 23957,
  27208, 27150, 26984, 26724, 26050, 24978, 23625, 22871, 22473, 22573, 
    22788, 23383, 24362, 25491, 26424, 27201, 26979, 26415, 26019, 25373, 
    24495, 23976,
  27089, 27066, 26832, 26675, 26075, 25020, 23684, 22883, 22484, 22556, 
    22891, 23413, 24221, 25509, 26431, 27045, 26835, 26394, 25950, 25448, 
    24609, 23876,
  26887, 26874, 26851, 26675, 26070, 25045, 23684, 22915, 22513, 22552, 
    22845, 23496, 24349, 25344, 26720, 26914, 26531, 26184, 25867, 25441, 
    24666, 24103,
  26634, 26599, 26771, 26592, 26070, 25076, 23743, 22959, 22545, 22564, 
    22867, 23445, 24263, 25261, 26429, 26889, 26513, 26134, 25776, 25404, 
    24748, 24103,
  26387, 26321, 26692, 26562, 26087, 25084, 23701, 22947, 22542, 22552, 
    22810, 23419, 24203, 25340, 26819, 26934, 26637, 26220, 25915, 25485, 
    24710, 24183,
  26203, 26133, 26694, 26572, 26113, 25143, 23816, 23009, 22618, 22626, 
    22890, 23414, 24351, 25412, 26510, 27021, 26854, 26393, 25984, 25534, 
    24824, 24216,
  26115, 26072, 26687, 26591, 26138, 25123, 23805, 22994, 22629, 22560, 
    22830, 23447, 24245, 25255, 26224, 27054, 26917, 26479, 26101, 25632, 
    24881, 24396,
  26110, 26093, 26610, 26610, 26154, 25103, 23791, 23023, 22562, 22623, 
    22801, 23482, 24237, 25344, 26712, 27093, 27048, 26551, 26114, 25670, 
    24976, 24283,
  26143, 26117, 26623, 26582, 26121, 25159, 23836, 23064, 22585, 22657, 
    22937, 23424, 24373, 25299, 26654, 27065, 27210, 26595, 26176, 25776, 
    25078, 24389,
  26165, 26093, 26575, 26556, 26143, 25181, 23871, 23076, 22620, 22585, 
    22797, 23482, 24146, 25472, 26372, 26885, 26823, 26443, 26162, 25657, 
    24950, 24463,
  26154, 26030, 26524, 26529, 26157, 25190, 23874, 23084, 22672, 22599, 
    22943, 23362, 24197, 25371, 26753, 26823, 26742, 26320, 25996, 25570, 
    24925, 24376,
  26115, 25962, 26451, 26572, 26151, 25235, 23884, 23081, 22672, 22613, 
    22908, 23436, 24241, 25139, 26697, 26840, 27197, 26616, 26259, 25819, 
    25141, 24549,
  26074, 25926, 26509, 26534, 26209, 25246, 23887, 23140, 22704, 22608, 
    22891, 23410, 24330, 25364, 26620, 26913, 27216, 26695, 26334, 25900, 
    25275, 24777,
  26080, 25959, 26514, 26529, 26146, 25279, 23925, 23155, 22715, 22642, 
    22802, 23499, 24286, 25201, 26107, 26866, 27110, 26651, 26299, 25874, 
    25300, 24891,
  26179, 26098, 26510, 26475, 26135, 25226, 23960, 23149, 22733, 22627, 
    22837, 23392, 24184, 25362, 26257, 26824, 27079, 26572, 26292, 25906, 
    25376, 24871,
  26378, 26346, 26684, 26540, 26106, 25187, 23932, 23169, 22721, 22581, 
    22865, 23400, 24280, 25257, 26500, 26888, 26879, 26370, 26175, 25843, 
    25421, 24951,
  26624, 26641, 26826, 26601, 26134, 25169, 23960, 23137, 22771, 22647, 
    22916, 23407, 24078, 25354, 26598, 26960, 26773, 26399, 26147, 25781, 
    25414, 25004,
  26835, 26887, 26864, 26650, 26172, 25172, 23932, 23166, 22741, 22647, 
    22788, 23417, 24272, 25487, 26563, 26963, 26710, 26326, 26057, 25613, 
    25338, 25011,
  26952, 27024, 26922, 26682, 26175, 25212, 23914, 23160, 22797, 22663, 
    22839, 23353, 24203, 25377, 26342, 26982, 26742, 26247, 25989, 25600, 
    25274, 24991,
  26978, 27067, 26970, 26735, 26172, 25220, 23942, 23186, 22717, 22689, 
    22938, 23363, 24169, 25091, 26439, 27035, 26748, 26225, 25913, 25557, 
    25101, 24903,
  26964, 27067, 27029, 26793, 26185, 25257, 23956, 23222, 22791, 22643, 
    22830, 23447, 24097, 25419, 26675, 27032, 26835, 26240, 25843, 25351, 
    25038, 24742,
  26962, 27065, 27029, 26810, 26209, 25242, 23987, 23207, 22761, 22686, 
    22921, 23434, 24102, 25366, 26371, 27017, 26879, 26254, 25843, 25426, 
    25025, 24695,
  26985, 27067, 27029, 26768, 26237, 25276, 24008, 23245, 22829, 22640, 
    22850, 23394, 24038, 25438, 26345, 27017, 26773, 26101, 25754, 25320, 
    24903, 24575,
  26998, 27054, 26937, 26825, 26282, 25262, 23990, 23195, 22823, 22695, 
    22898, 23442, 24178, 25382, 26760, 26954, 26742, 26023, 25609, 25282, 
    24859, 24494,
  26967, 27007, 27003, 26822, 26294, 25265, 24008, 23221, 22802, 22712, 
    22833, 23348, 24181, 25168, 26534, 26916, 25925, 25424, 25298, 25002, 
    24610, 24313,
  26880, 26917, 26973, 26798, 26300, 25284, 24022, 23233, 22810, 22654, 
    22832, 23368, 24159, 25382, 26298, 26794, 25377, 24954, 24904, 24828, 
    24470, 24192,
  26720, 26769, 27003, 26832, 26282, 25332, 23980, 23254, 22761, 22706, 
    22847, 23373, 24230, 25329, 26456, 26829, 25595, 25149, 24994, 24766, 
    24476, 24125,
  26453, 26524, 26942, 26787, 26263, 25270, 23987, 23251, 22825, 22712, 
    22915, 23330, 24163, 25347, 26293, 26851, 26324, 25734, 25484, 24996, 
    24572, 24192,
  26076, 26167, 26656, 26579, 26207, 25309, 24004, 23251, 22834, 22697, 
    22880, 23345, 24237, 25312, 26609, 26601, 25987, 25423, 25139, 24871, 
    24534, 24212,
  25668, 25760, 26346, 26404, 26062, 25265, 23973, 23257, 22773, 22760, 
    22887, 23426, 24282, 25259, 26347, 26248, 25832, 25409, 25180, 24772, 
    24515, 24118,
  25355, 25430, 26176, 26316, 26045, 25247, 23990, 23254, 22852, 22792, 
    22992, 23411, 24193, 25333, 26676, 26087, 26374, 25828, 25491, 25058, 
    24585, 24131,
  25238, 25293, 26143, 26301, 26031, 25211, 23986, 23227, 22840, 22734, 
    22921, 23342, 24133, 25493, 26568, 26009, 26748, 26332, 25863, 25400, 
    24776, 24266,
  25329, 25380, 26132, 26275, 26082, 25267, 23973, 23268, 22804, 22798, 
    22898, 23386, 24129, 25249, 26801, 26014, 26760, 26535, 26050, 25475, 
    24820, 24393,
  25555, 25620, 26368, 26407, 26145, 25267, 23993, 23254, 22831, 22749, 
    22880, 23401, 24089, 25375, 26560, 26393, 26972, 26635, 26104, 25575, 
    24916, 24353,
  25790, 25872, 26688, 26651, 26266, 25287, 23976, 23242, 22799, 22789, 
    22929, 23431, 24062, 25224, 26298, 26829, 27365, 26810, 26209, 25631, 
    24865, 24393,
  25912, 25994, 26874, 26719, 26300, 25298, 23990, 23239, 22837, 22737, 
    22983, 23436, 24245, 25323, 26310, 26994, 27482, 26774, 26209, 25654, 
    24929, 24454,
  25837, 25909, 26737, 26647, 26197, 25281, 23983, 23251, 22875, 22726, 
    22898, 23386, 24358, 25287, 26726, 26882, 27365, 26831, 26278, 25754, 
    24916, 24447,
  25527, 25605, 26534, 26501, 26140, 25281, 23983, 23277, 22855, 22706, 
    23020, 23373, 24190, 25251, 26504, 26638, 27201, 26860, 26320, 25774, 
    25101, 24588,
  24964, 25078, 26363, 26445, 26117, 25217, 23963, 23239, 22866, 22798, 
    22924, 23399, 24289, 25329, 26369, 26479, 27221, 26875, 26396, 25824, 
    25095, 24474,
  24155, 24328, 26098, 26216, 26004, 25209, 23945, 23227, 22858, 22726, 
    22869, 23302, 24287, 25375, 26551, 26309, 27172, 26853, 26354, 25829, 
    25107, 24554,
  23157, 23397, 25635, 25954, 25831, 25093, 23924, 23198, 22867, 22789, 
    22910, 23363, 24095, 25352, 25926, 25829, 27041, 26751, 26360, 25756, 
    25082, 24447,
  22105, 22408, 24718, 25319, 25590, 25032, 23900, 23234, 22858, 22775, 
    22915, 23422, 24216, 25331, 26619, 24778, 26585, 26679, 26326, 25818, 
    25101, 24387,
  21196, 21535, 23903, 24788, 25384, 24996, 23907, 23219, 22820, 22819, 
    22870, 23473, 24161, 25212, 26214, 23705, 25782, 26564, 26285, 25779, 
    25057, 24568,
  20614, 20947, 23612, 24594, 25267, 24956, 23897, 23249, 22849, 22847, 
    23010, 23336, 24290, 25273, 26340, 23277, 25714, 26522, 26320, 25868, 
    25217, 24608,
  20458, 20755, 23807, 24643, 25279, 24894, 23894, 23237, 22897, 22798, 
    22998, 23455, 24223, 25243, 26449, 23279, 25645, 26594, 26360, 25918, 
    25261, 24622,
  20700, 20956, 23916, 24778, 25318, 24951, 23870, 23202, 22850, 22782, 
    22944, 23471, 24243, 25499, 26532, 23669, 25832, 26615, 26410, 25879, 
    25242, 24723,
  21197, 21403, 24183, 24939, 25367, 24872, 23870, 23181, 22832, 22825, 
    23016, 23371, 24007, 25319, 26471, 23986, 25920, 26572, 26341, 25918, 
    25319, 24823,
  21736, 21879, 24447, 25080, 25399, 24915, 23852, 23190, 22853, 22810, 
    23025, 23412, 24293, 25431, 26573, 24231, 25988, 26594, 26314, 25929, 
    25325, 24743,
  22134, 22227, 24457, 25118, 25339, 24859, 23811, 23155, 22850, 22877, 
    23002, 23451, 24308, 25550, 26124, 24194, 25851, 26515, 26326, 25843, 
    25217, 24683,
  22325, 22407, 24368, 25085, 25334, 24859, 23825, 23182, 22865, 22854, 
    23053, 23466, 24246, 25606, 26591, 24060, 25732, 26443, 26238, 25806, 
    25236, 24710,
  22356, 22449, 24371, 25023, 25296, 24808, 23804, 23143, 22839, 22814, 
    22980, 23444, 24350, 25378, 26345, 24040, 25845, 26421, 26182, 25713, 
    25129, 24697,
  22291, 22375, 24333, 25056, 25328, 24758, 23738, 23123, 22827, 22877, 
    23082, 23502, 24330, 25429, 26384, 24048, 25757, 26500, 26217, 25788, 
    25109, 24630,
  22134, 22191, 24457, 25085, 25308, 24806, 23710, 23129, 22886, 22837, 
    23156, 23408, 24427, 25272, 26913, 24299, 26007, 26443, 26217, 25689, 
    25231, 24831,
  21855, 21908, 24338, 25040, 25282, 24786, 23721, 23171, 22898, 22809, 
    23080, 23459, 24378, 25574, 26737, 24401, 26144, 26537, 26231, 25732, 
    25199, 24805,
  21481, 21575, 23991, 24787, 25197, 24711, 23704, 23180, 22898, 22858, 
    23095, 23548, 24316, 25409, 26297, 23994, 25957, 26494, 26176, 25770, 
    25244, 24772,
  21138, 21288, 23646, 24596, 25162, 24750, 23732, 23189, 22901, 22852, 
    23009, 23599, 24237, 25520, 26503, 23627, 25671, 26479, 26210, 25701, 
    25314, 24832,
  20984, 21158, 23639, 24642, 25154, 24714, 23704, 23162, 22887, 22919, 
    22995, 23592, 24393, 25369, 26807, 23629, 25796, 26335, 26107, 25751, 
    25206, 24745,
  21082, 21244, 23966, 24765, 25194, 24675, 23687, 23195, 22905, 22936, 
    23124, 23600, 24364, 25583, 26545, 23896, 25926, 26307, 26101, 25707, 
    25219, 24705,
  21336, 21500, 24265, 24960, 25223, 24680, 23663, 23154, 22911, 22950, 
    23067, 23577, 24423, 25500, 26938, 24319, 26039, 26379, 26129, 25640, 
    25079, 24632,
  21564, 21780, 24555, 25084, 25214, 24627, 23635, 23136, 22911, 22965, 
    23081, 23547, 24393, 25642, 26582, 24611, 26232, 26335, 26046, 25572, 
    25118, 24699,
  21636, 21929, 24560, 25135, 25240, 24602, 23646, 23116, 22949, 22968, 
    23099, 23631, 24436, 25757, 26785, 24603, 26164, 26329, 26019, 25622, 
    24991, 24612,
  21556, 21888, 24499, 25133, 25252, 24597, 23618, 23113, 22941, 22980, 
    23087, 23494, 24510, 25668, 27409, 24427, 26082, 26329, 26004, 25560, 
    25023, 24465,
  21436, 21735, 24484, 25092, 25212, 24594, 23588, 23137, 22947, 22946, 
    23051, 23591, 24444, 25721, 26909, 24278, 26015, 26335, 25978, 25517, 
    24921, 24512,
  21409, 21625, 24522, 25084, 25180, 24522, 23546, 23094, 22915, 22926, 
    23014, 23639, 24542, 25726, 27021, 24214, 25940, 26322, 25999, 25617, 
    24947, 24506,
  21540, 21667, 24525, 25092, 25195, 24497, 23526, 23079, 22947, 22975, 
    23222, 23634, 24693, 25845, 26810, 24138, 25872, 26315, 26075, 25573, 
    25126, 24693,
  21809, 21870, 24571, 25149, 25149, 24458, 23505, 23138, 22942, 22998, 
    23140, 23619, 24459, 25889, 26701, 24077, 25922, 26337, 26054, 25698, 
    25120, 24661,
  22145, 22172, 24635, 25187, 25132, 24418, 23467, 23085, 22939, 23047, 
    23126, 23653, 24511, 25787, 26807, 24163, 25898, 26235, 26034, 25610, 
    25120, 24694,
  22471, 22495, 24779, 25198, 25141, 24396, 23460, 23068, 22933, 23007, 
    23194, 23678, 24486, 25668, 27031, 24268, 25916, 26316, 26013, 25692, 
    25139, 24728,
  22748, 22783, 24838, 25241, 25147, 24352, 23474, 23098, 22934, 23022, 
    23283, 23645, 24519, 25851, 26716, 24307, 25947, 26279, 25993, 25660, 
    25082, 24541,
  22983, 23023, 24932, 25295, 25107, 24310, 23429, 23057, 22995, 23025, 
    23098, 23793, 24548, 25845, 27121, 24371, 25979, 26229, 25917, 25580, 
    25133, 24581,
  23209, 23243, 25069, 25338, 25104, 24268, 23423, 23080, 22978, 23026, 
    23209, 23712, 24465, 25718, 27035, 24451, 26054, 26179, 25924, 25562, 
    25006, 24521,
  23448, 23463, 25190, 25414, 25053, 24246, 23406, 23104, 22949, 22989, 
    23181, 23657, 24611, 25839, 27035, 24479, 26072, 26207, 25869, 25450, 
    24930, 24502,
  23707, 23683, 25307, 25398, 25044, 24139, 23367, 23054, 22976, 23035, 
    23184, 23695, 24621, 25825, 26876, 24548, 26016, 26173, 25849, 25451, 
    24988, 24448,
  23994, 23917, 25373, 25360, 24985, 24123, 23319, 23096, 23011, 23015, 
    23224, 23789, 24707, 25837, 26571, 24503, 25954, 26122, 25774, 25383, 
    24867, 24375,
  24276, 24159, 25348, 25406, 24942, 24064, 23267, 23061, 22997, 23061, 
    23188, 23795, 24692, 25982, 26957, 24539, 25967, 26057, 25684, 25364, 
    24836, 24282,
  24420, 24298, 25386, 25347, 24845, 24017, 23268, 23082, 22968, 23007, 
    23208, 23825, 24639, 25829, 26932, 24634, 25974, 25928, 25616, 25303, 
    24709, 24222,
  24299, 24190, 25452, 25382, 24771, 23913, 23240, 23002, 22994, 23018, 
    23177, 23881, 24703, 26046, 27241, 24756, 25968, 25813, 25540, 25172, 
    24601, 24055,
  24008, 23903, 25447, 25310, 24739, 23916, 23206, 23041, 22989, 23013, 
    23234, 23864, 24885, 26118, 27110, 24862, 26079, 25770, 25430, 25024, 
    24494, 23962,
  23853, 23746, 25462, 25286, 24708, 23841, 23165, 23044, 22972, 23139, 
    23243, 23882, 24876, 26141, 27350, 24800, 26085, 25734, 25313, 24881, 
    24322, 23815,
  27970, 27902, 27257, 26693, 25583, 24079, 22720, 22262, 22193, 22516, 
    22864, 23671, 24671, 25882, 26493, 27735, 27140, 26226, 25679, 25031, 
    24187, 23592,
  27916, 27844, 27134, 26682, 25623, 24185, 22820, 22256, 22166, 22556, 
    22853, 23590, 24578, 25543, 26835, 27572, 26978, 26024, 25534, 25043, 
    24378, 23805,
  27801, 27726, 27040, 26537, 25591, 24249, 22914, 22303, 22180, 22507, 
    22835, 23592, 24587, 25399, 26593, 27225, 26816, 26081, 25657, 25111, 
    24454, 23918,
  27702, 27643, 26900, 26467, 25637, 24319, 22948, 22382, 22236, 22512, 
    22886, 23660, 24560, 25651, 26634, 26966, 26654, 26125, 25734, 25192, 
    24555, 23905,
  27642, 27612, 26771, 26442, 25634, 24394, 23017, 22411, 22221, 22446, 
    22948, 23634, 24609, 25847, 26910, 26667, 26299, 25887, 25568, 25185, 
    24491, 23945,
  27605, 27581, 26710, 26418, 25637, 24425, 23097, 22458, 22255, 22506, 
    22909, 23523, 24515, 25738, 26823, 26379, 25117, 25123, 25141, 24924, 
    24376, 23924,
  27576, 27521, 26799, 26493, 25742, 24512, 23138, 22543, 22273, 22560, 
    22879, 23594, 24574, 25851, 26535, 26489, 25440, 25396, 25216, 24918, 
    24433, 23871,
  27541, 27448, 26981, 26609, 25840, 24590, 23211, 22587, 22255, 22525, 
    22871, 23560, 24448, 25628, 26701, 26794, 25957, 25569, 25347, 24898, 
    24357, 23937,
  27477, 27384, 27073, 26726, 25907, 24730, 23283, 22578, 22340, 22542, 
    22862, 23520, 24416, 25607, 26794, 27095, 26598, 25907, 25512, 24948, 
    24382, 23870,
  27374, 27316, 27110, 26732, 25976, 24738, 23315, 22657, 22348, 22459, 
    22853, 23577, 24440, 25723, 26587, 27343, 26996, 26095, 25491, 24948, 
    24311, 23796,
  27245, 27226, 27044, 26762, 26007, 24797, 23345, 22671, 22315, 22479, 
    22847, 23437, 24497, 25393, 26774, 27374, 26871, 25979, 25456, 24854, 
    24260, 23822,
  27114, 27126, 27001, 26726, 25962, 24802, 23418, 22721, 22377, 22573, 
    22801, 23524, 24381, 25674, 26766, 27316, 26771, 25914, 25456, 24916, 
    24374, 23882,
  27017, 27045, 26996, 26689, 26016, 24833, 23435, 22733, 22388, 22570, 
    22790, 23529, 24329, 25500, 26254, 27271, 26815, 26123, 25566, 24978, 
    24380, 23868,
  26988, 27008, 26900, 26635, 25993, 24866, 23515, 22730, 22420, 22578, 
    22898, 23450, 24287, 25660, 26412, 27263, 27064, 26281, 25766, 25226, 
    24539, 23988,
  27032, 27022, 26943, 26676, 26087, 24925, 23546, 22797, 22400, 22483, 
    22840, 23505, 24402, 25601, 26496, 27279, 27257, 26510, 26007, 25319, 
    24469, 24022,
  27112, 27069, 26993, 26732, 26096, 24953, 23566, 22821, 22425, 22552, 
    22877, 23477, 24281, 25551, 26310, 27289, 27170, 26504, 25985, 25356, 
    24577, 23914,
  27169, 27117, 27010, 26772, 26070, 24989, 23594, 22802, 22422, 22517, 
    22752, 23484, 24306, 25531, 26562, 27229, 26871, 26418, 25985, 25380, 
    24614, 23974,
  27156, 27126, 26929, 26718, 26060, 25011, 23639, 22891, 22457, 22545, 
    22794, 23400, 24387, 25429, 26467, 27116, 26901, 26410, 25923, 25399, 
    24538, 24027,
  27052, 27046, 26892, 26659, 26057, 24989, 23653, 22885, 22518, 22548, 
    22825, 23415, 24381, 25566, 26607, 26988, 26696, 26279, 25923, 25430, 
    24710, 24087,
  26859, 26852, 26734, 26592, 26090, 25014, 23656, 22940, 22462, 22536, 
    22850, 23420, 24211, 25471, 26560, 26910, 26322, 26135, 25903, 25442, 
    24684, 24087,
  26616, 26582, 26722, 26594, 26035, 25062, 23718, 22958, 22588, 22556, 
    22862, 23405, 24332, 25401, 26637, 26921, 26609, 26316, 26006, 25529, 
    24849, 24160,
  26387, 26323, 26656, 26538, 26087, 25075, 23746, 22973, 22547, 22567, 
    22853, 23371, 24184, 25189, 26348, 26985, 26676, 26345, 25971, 25504, 
    24893, 24180,
  26233, 26165, 26617, 26482, 26107, 25100, 23749, 22978, 22573, 22567, 
    22927, 23463, 24294, 25345, 26391, 26985, 26832, 26344, 26040, 25584, 
    24861, 24240,
  26178, 26134, 26574, 26551, 26112, 25117, 23790, 23028, 22570, 22618, 
    22858, 23406, 24309, 25484, 26173, 27025, 26882, 26453, 26116, 25609, 
    24886, 24320,
  26192, 26178, 26622, 26548, 26124, 25139, 23794, 23016, 22628, 22600, 
    22866, 23409, 24262, 25312, 26488, 27003, 26976, 26525, 26226, 25751, 
    25071, 24421,
  26220, 26207, 26635, 26589, 26115, 25139, 23825, 23086, 22616, 22566, 
    22838, 23429, 24375, 25547, 26639, 26950, 27082, 26610, 26253, 25826, 
    25090, 24541,
  26219, 26166, 26632, 26594, 26121, 25153, 23874, 23083, 22607, 22612, 
    22818, 23367, 24227, 25251, 26557, 26785, 26451, 26272, 26046, 25707, 
    25045, 24621,
  26172, 26064, 26637, 26569, 26101, 25209, 23898, 23104, 22677, 22634, 
    22863, 23406, 24271, 25460, 26471, 26826, 26788, 26379, 26122, 25689, 
    25128, 24540,
  26094, 25950, 26566, 26518, 26121, 25195, 23873, 23101, 22636, 22591, 
    22854, 23410, 24266, 25419, 26459, 26892, 27287, 26719, 26307, 25838, 
    25204, 24735,
  26020, 25876, 26518, 26501, 26115, 25242, 23859, 23130, 22650, 22597, 
    22860, 23293, 24118, 25419, 26713, 26914, 27249, 26639, 26253, 25857, 
    25268, 24788,
  26003, 25886, 26419, 26434, 26129, 25192, 23855, 23095, 22674, 22625, 
    22894, 23316, 24083, 25265, 26779, 26803, 27106, 26603, 26266, 25857, 
    25408, 24862,
  26097, 26024, 26451, 26415, 26100, 25183, 23894, 23118, 22715, 22590, 
    22805, 23446, 24127, 25255, 26360, 26707, 27062, 26545, 26190, 25869, 
    25464, 25117,
  26324, 26298, 26557, 26515, 26034, 25172, 23880, 23109, 22712, 22651, 
    22950, 23453, 24224, 25339, 26242, 26800, 26832, 26379, 26149, 25838, 
    25439, 25123,
  26639, 26653, 26789, 26688, 26151, 25236, 23939, 23129, 22755, 22677, 
    22819, 23448, 24150, 25344, 26126, 26925, 26744, 26278, 26010, 25701, 
    25343, 24995,
  26946, 26986, 26964, 26706, 26166, 25155, 23928, 23159, 22761, 22642, 
    22850, 23328, 24105, 25425, 26587, 26962, 26694, 26235, 25976, 25663, 
    25343, 24901,
  27157, 27220, 26942, 26771, 26185, 25197, 23921, 23161, 22720, 22691, 
    22899, 23379, 24127, 25330, 26490, 26973, 26626, 26132, 25865, 25483, 
    25171, 24928,
  27247, 27343, 27038, 26793, 26217, 25222, 23914, 23215, 22804, 22653, 
    22870, 23330, 24092, 25362, 26706, 26917, 25978, 25599, 25396, 25177, 
    24795, 24478,
  27261, 27389, 27023, 26763, 26192, 25244, 23949, 23214, 22758, 22710, 
    22864, 23427, 24174, 25330, 26332, 26965, 26021, 25526, 25292, 25009, 
    24635, 24371,
  27257, 27390, 26967, 26814, 26237, 25247, 23969, 23226, 22784, 22610, 
    22841, 23355, 24324, 25185, 26535, 26951, 26582, 25873, 25548, 25165, 
    24743, 24371,
  27251, 27353, 27007, 26776, 26226, 25281, 23973, 23214, 22822, 22704, 
    22898, 23345, 24142, 25243, 26670, 26909, 26432, 25866, 25582, 25271, 
    24794, 24499,
  27209, 27263, 26907, 26757, 26220, 25259, 23976, 23211, 22807, 22704, 
    22989, 23370, 24260, 25441, 26815, 26856, 25921, 25541, 25258, 25102, 
    24679, 24351,
  27081, 27100, 26959, 26787, 26246, 25267, 23986, 23241, 22828, 22693, 
    22872, 23261, 24211, 25387, 25994, 26842, 25909, 25411, 25195, 24897, 
    24629, 24243,
  26841, 26850, 26944, 26728, 26237, 25286, 23979, 23217, 22769, 22658, 
    22952, 23312, 24028, 25350, 26419, 26859, 26675, 25951, 25637, 25183, 
    24749, 24297,
  26484, 26505, 26771, 26741, 26234, 25284, 23979, 23253, 22825, 22690, 
    22895, 23431, 24181, 25194, 26793, 26884, 26706, 26053, 25664, 25258, 
    24692, 24451,
  26017, 26069, 26651, 26609, 26206, 25303, 24004, 23273, 22813, 22750, 
    22995, 23421, 24213, 25266, 26796, 26706, 26725, 26075, 25623, 25171, 
    24673, 24384,
  25493, 25573, 26354, 26453, 26137, 25236, 23976, 23226, 22851, 22698, 
    22887, 23398, 24230, 25250, 26446, 26389, 26582, 25995, 25575, 25208, 
    24622, 24290,
  25017, 25106, 26051, 26243, 26010, 25216, 24028, 23294, 22851, 22724, 
    22926, 23281, 24267, 25241, 26468, 26054, 26438, 26191, 25664, 25196, 
    24654, 24297,
  24710, 24784, 25914, 26194, 26054, 25230, 24018, 23241, 22854, 22776, 
    22938, 23396, 24213, 25087, 26412, 25882, 26806, 26414, 25920, 25295, 
    24769, 24250,
  24630, 24682, 25901, 26194, 26034, 25272, 23983, 23309, 22813, 22710, 
    22938, 23426, 24119, 25245, 26672, 25849, 26937, 26696, 26141, 25519, 
    24845, 24391,
  24744, 24794, 26114, 26299, 26082, 25267, 24011, 23250, 22851, 22681, 
    22858, 23462, 24247, 25339, 26407, 26018, 27162, 26790, 26189, 25675, 
    24928, 24484,
  24947, 25022, 26340, 26396, 26179, 25264, 23959, 23235, 22825, 22732, 
    22880, 23376, 24154, 25217, 26397, 26357, 27229, 26804, 26265, 25656, 
    25011, 24471,
  25114, 25216, 26441, 26472, 26137, 25278, 23997, 23276, 22825, 22776, 
    22943, 23482, 24166, 25257, 26579, 26517, 27274, 26775, 26257, 25637, 
    24972, 24444,
  25143, 25244, 26528, 26531, 26197, 25227, 23969, 23238, 22865, 22779, 
    22921, 23320, 24284, 25481, 26315, 26667, 27285, 26782, 26285, 25712, 
    25017, 24464,
  24975, 25059, 26548, 26542, 26171, 25255, 23972, 23285, 22866, 22787, 
    22943, 23363, 24230, 25408, 26473, 26756, 27385, 26848, 26300, 25700, 
    24985, 24431,
  24597, 24685, 26398, 26372, 26145, 25261, 23955, 23211, 22845, 22776, 
    22929, 23439, 24252, 25527, 26720, 26553, 27379, 26768, 26307, 25731, 
    25023, 24425,
  24026, 24157, 25987, 26156, 25939, 25149, 23945, 23276, 22871, 22710, 
    22949, 23465, 24124, 25215, 26479, 26213, 27193, 26819, 26259, 25781, 
    25062, 24438,
  23303, 23495, 25528, 25787, 25828, 25118, 23938, 23241, 22883, 22736, 
    22858, 23381, 24171, 25264, 26839, 25818, 27012, 26760, 26265, 25775, 
    25170, 24499,
  22504, 22745, 24986, 25442, 25639, 25082, 23927, 23262, 22837, 22848, 
    22930, 23379, 24274, 25315, 26300, 25166, 26644, 26682, 26259, 25825, 
    25069, 24552,
  21742, 22013, 24174, 24971, 25396, 24989, 23927, 23288, 22860, 22773, 
    22967, 23437, 24265, 25360, 26597, 24214, 25953, 26581, 26231, 25800, 
    25050, 24586,
  21156, 21432, 23872, 24702, 25315, 24990, 23883, 23259, 22869, 22771, 
    22984, 23381, 24196, 25430, 26510, 23623, 25710, 26581, 26300, 25887, 
    25222, 24539,
  20860, 21115, 23979, 24815, 25356, 24990, 23900, 23223, 22860, 22785, 
    22953, 23488, 24231, 25206, 26531, 23673, 25878, 26551, 26335, 25887, 
    25164, 24646,
  20889, 21116, 24204, 24934, 25353, 24936, 23907, 23229, 22905, 22797, 
    23021, 23336, 24253, 25306, 26490, 23988, 26028, 26596, 26328, 25837, 
    25164, 24693,
  21187, 21396, 24275, 24947, 25362, 24922, 23844, 23200, 22872, 22782, 
    23021, 23463, 24154, 25299, 26898, 24093, 26090, 26559, 26251, 25868, 
    25171, 24626,
  21632, 21818, 24299, 24988, 25353, 24934, 23841, 23195, 22890, 22817, 
    22962, 23481, 24263, 25325, 26404, 24076, 25741, 26531, 26266, 25850, 
    25241, 24734,
  22073, 22210, 24514, 25090, 25405, 24883, 23848, 23189, 22855, 22803, 
    23022, 23430, 24160, 25355, 26750, 24215, 25854, 26603, 26294, 25838, 
    25171, 24721,
  22384, 22474, 24611, 25139, 25411, 24850, 23838, 23159, 22864, 22789, 
    22945, 23458, 24224, 25453, 26600, 24301, 25804, 26582, 26253, 25800, 
    25184, 24667,
  22521, 22603, 24593, 25157, 25387, 24864, 23797, 23201, 22917, 22883, 
    23022, 23420, 24234, 25421, 26592, 24218, 25791, 26466, 26197, 25794, 
    25159, 24701,
  22519, 22617, 24507, 25109, 25376, 24861, 23814, 23154, 22908, 22838, 
    22988, 23461, 24296, 25402, 27020, 24122, 25767, 26466, 26225, 25738, 
    25121, 24634,
  22418, 22514, 24421, 25080, 25385, 24836, 23807, 23213, 22912, 22832, 
    22945, 23428, 24298, 25538, 26593, 24081, 25854, 26429, 26218, 25751, 
    25147, 24681,
  22205, 22280, 24444, 25144, 25402, 24819, 23759, 23169, 22868, 22887, 
    23017, 23433, 24385, 25591, 26549, 24347, 26047, 26517, 26218, 25696, 
    25122, 24755,
  21857, 21927, 24310, 25021, 25334, 24760, 23731, 23184, 22929, 22864, 
    22949, 23515, 24254, 25480, 26884, 24297, 25967, 26429, 26198, 25739, 
    25109, 24782,
  21416, 21518, 23914, 24781, 25225, 24749, 23703, 23178, 22871, 22836, 
    23080, 23523, 24397, 25377, 26532, 23868, 25785, 26467, 26143, 25746, 
    25185, 24716,
  21031, 21179, 23669, 24689, 25134, 24671, 23673, 23140, 22927, 22870, 
    23055, 23432, 24316, 25403, 26644, 23511, 25668, 26316, 26053, 25651, 
    25192, 24629,
  20875, 21042, 23752, 24660, 25148, 24671, 23690, 23126, 22898, 22868, 
    23018, 23495, 24393, 25600, 26707, 23608, 25785, 26323, 25971, 25497, 
    24995, 24622,
  21017, 21170, 23975, 24792, 25154, 24722, 23697, 23167, 22901, 22874, 
    23038, 23534, 24226, 25468, 26560, 23886, 25873, 26294, 25950, 25560, 
    24969, 24562,
  21357, 21504, 24173, 24946, 25223, 24683, 23659, 23152, 22966, 22909, 
    23072, 23618, 24452, 25789, 26960, 24240, 25973, 26374, 26068, 25603, 
    24989, 24435,
  21708, 21891, 24437, 25035, 25254, 24607, 23625, 23121, 22945, 22895, 
    23081, 23674, 24367, 25731, 26887, 24504, 26067, 26323, 26006, 25560, 
    25008, 24556,
  21926, 22170, 24569, 25140, 25234, 24616, 23594, 23127, 22943, 22895, 
    23161, 23532, 24381, 25550, 27084, 24601, 26148, 26381, 26041, 25629, 
    24983, 24469,
  21984, 22267, 24681, 25170, 25240, 24551, 23625, 23142, 22949, 22924, 
    23201, 23659, 24350, 25682, 26892, 24646, 26148, 26287, 26041, 25579, 
    24926, 24436,
  21960, 22233, 24693, 25164, 25218, 24554, 23580, 23124, 22920, 22932, 
    23076, 23588, 24370, 25583, 26890, 24542, 26060, 26317, 26000, 25561, 
    25028, 24557,
  21954, 22184, 24686, 25183, 25223, 24518, 23532, 23139, 22888, 22956, 
    23060, 23596, 24375, 25676, 26882, 24433, 25974, 26324, 25951, 25629, 
    24991, 24470,
  22024, 22204, 24661, 25154, 25183, 24482, 23497, 23116, 22970, 22941, 
    23145, 23660, 24459, 25818, 26846, 24279, 25949, 26301, 26069, 25717, 
    25188, 24524,
  22165, 22296, 24641, 25152, 25172, 24468, 23511, 23089, 22979, 22942, 
    23060, 23617, 24434, 25937, 26851, 24234, 25856, 26295, 26021, 25679, 
    25156, 24531,
  22341, 22431, 24679, 25141, 25144, 24398, 23477, 23125, 22974, 22957, 
    23203, 23561, 24612, 25718, 26760, 24178, 25856, 26296, 26042, 25717, 
    25112, 24665,
  22526, 22589, 24748, 25168, 25144, 24376, 23470, 23096, 22924, 22977, 
    23103, 23587, 24592, 25684, 26817, 24211, 25881, 26238, 25973, 25649, 
    25055, 24652,
  22719, 22766, 24809, 25230, 25147, 24345, 23457, 23084, 23000, 23035, 
    23024, 23691, 24640, 25516, 26616, 24325, 26037, 26318, 25987, 25606, 
    24992, 24404,
  22940, 22971, 24979, 25327, 25110, 24334, 23460, 23076, 23021, 23020, 
    23158, 23608, 24581, 25737, 27009, 24434, 26056, 26231, 25960, 25531, 
    24948, 24519,
  23204, 23213, 25103, 25378, 25122, 24304, 23436, 23091, 22983, 23049, 
    23167, 23643, 24551, 25749, 26699, 24544, 26187, 26203, 25904, 25637, 
    25056, 24499,
  23495, 23483, 25245, 25446, 25016, 24245, 23398, 23091, 22975, 22989, 
    23181, 23735, 24670, 25728, 26876, 24692, 26156, 26138, 25898, 25538, 
    25012, 24405,
  23788, 23752, 25354, 25430, 25036, 24209, 23350, 23088, 22993, 23007, 
    23218, 23768, 24641, 25960, 27457, 24667, 26050, 26138, 25835, 25458, 
    24897, 24352,
  24080, 24007, 25418, 25403, 24965, 24139, 23322, 23074, 23051, 23039, 
    23222, 23769, 24744, 25928, 26979, 24518, 25976, 26038, 25692, 25328, 
    24809, 24232,
  24347, 24235, 25398, 25382, 24908, 24064, 23298, 23089, 23031, 23019, 
    23268, 23820, 24656, 25994, 26904, 24421, 25932, 26016, 25601, 25266, 
    24694, 24166,
  24476, 24343, 25461, 25371, 24865, 24047, 23267, 23060, 23002, 22985, 
    23290, 23825, 24924, 26035, 27196, 24493, 25851, 25916, 25631, 25223, 
    24657, 24179,
  24352, 24223, 25441, 25374, 24836, 23966, 23268, 23072, 23049, 23091, 
    23243, 23823, 24767, 26164, 27010, 24581, 25964, 25851, 25548, 25130, 
    24619, 24073,
  24067, 23951, 25489, 25309, 24737, 23880, 23237, 23081, 23032, 23046, 
    23217, 23808, 24802, 25929, 27124, 24695, 26045, 25785, 25418, 25000, 
    24479, 23959,
  23916, 23805, 25421, 25280, 24694, 23821, 23209, 23019, 22965, 23014, 
    23217, 23892, 24954, 26201, 26937, 24712, 26144, 25743, 25369, 24919, 
    24308, 23866,
  27914, 27863, 27163, 26637, 25566, 24073, 22729, 22262, 22203, 22520, 
    22886, 23663, 24687, 25915, 26851, 27635, 26906, 26003, 25406, 24934, 
    24152, 23661,
  27863, 27807, 27200, 26654, 25635, 24219, 22861, 22306, 22223, 22532, 
    22865, 23639, 24610, 25722, 26642, 27550, 26968, 25982, 25453, 24872, 
    24278, 23741,
  27755, 27695, 26976, 26507, 25563, 24266, 22892, 22329, 22199, 22457, 
    22922, 23634, 24502, 25688, 26703, 27220, 26763, 26017, 25564, 24971, 
    24310, 23647,
  27669, 27618, 26782, 26397, 25580, 24325, 22971, 22370, 22245, 22474, 
    22930, 23543, 24447, 25878, 26497, 26818, 26439, 26010, 25577, 25058, 
    24399, 23821,
  27631, 27596, 26734, 26349, 25563, 24333, 23044, 22397, 22242, 22551, 
    22973, 23525, 24462, 25534, 26671, 26489, 25673, 25505, 25281, 24859, 
    24233, 23619,
  27615, 27579, 26714, 26367, 25651, 24445, 23089, 22493, 22227, 22459, 
    22870, 23522, 24496, 25578, 26266, 26478, 24989, 25101, 25060, 24840, 
    24214, 23820,
  27597, 27543, 26929, 26576, 25791, 24486, 23130, 22502, 22274, 22519, 
    22875, 23509, 24363, 25580, 26707, 26838, 26226, 25707, 25356, 24908, 
    24334, 23719,
  27560, 27504, 27096, 26726, 25912, 24612, 23227, 22540, 22282, 22504, 
    22872, 23529, 24431, 25632, 26872, 27254, 26918, 26009, 25473, 24889, 
    24251, 23672,
  27498, 27470, 27129, 26814, 25957, 24702, 23251, 22637, 22320, 22544, 
    22852, 23450, 24537, 25617, 26518, 27445, 27010, 26031, 25404, 24870, 
    24200, 23638,
  27409, 27415, 27200, 26812, 26032, 24716, 23320, 22622, 22340, 22518, 
    22823, 23419, 24350, 25545, 26319, 27523, 27010, 25966, 25424, 24832, 
    24168, 23598,
  27298, 27325, 27129, 26795, 26040, 24772, 23369, 22695, 22369, 22549, 
    22851, 23495, 24396, 25698, 26896, 27484, 26879, 25821, 25299, 24732, 
    24174, 23684,
  27171, 27215, 27078, 26731, 26014, 24808, 23396, 22680, 22360, 22529, 
    22922, 23510, 24408, 25679, 26493, 27431, 26824, 25987, 25396, 24825, 
    24186, 23710,
  27054, 27115, 26994, 26703, 25976, 24844, 23420, 22733, 22413, 22528, 
    22840, 23513, 24378, 25532, 26789, 27307, 26929, 26189, 25664, 25005, 
    24313, 23857,
  26989, 27046, 26879, 26701, 26071, 24909, 23476, 22771, 22398, 22500, 
    22885, 23548, 24395, 25412, 26534, 27339, 27160, 26390, 25829, 25185, 
    24389, 23897,
  26998, 27019, 26931, 26671, 26074, 24956, 23496, 22791, 22461, 22522, 
    22833, 23435, 24272, 25460, 26426, 27320, 27253, 26592, 26064, 25340, 
    24484, 23857,
  27055, 27036, 26979, 26695, 26037, 24894, 23562, 22832, 22435, 22502, 
    22870, 23377, 24378, 25583, 26522, 27295, 27116, 26513, 26043, 25409, 
    24497, 23836,
  27108, 27074, 26946, 26725, 26054, 24933, 23600, 22820, 22464, 22496, 
    22847, 23410, 24348, 25346, 26679, 27217, 27004, 26397, 25953, 25309, 
    24528, 23876,
  27110, 27081, 26997, 26710, 26056, 24983, 23641, 22858, 22502, 22553, 
    22849, 23399, 24407, 25476, 26682, 27169, 27004, 26353, 25918, 25302, 
    24496, 23929,
  27030, 27003, 26829, 26700, 26056, 24974, 23638, 22870, 22519, 22544, 
    22838, 23524, 24301, 25462, 26619, 27075, 26942, 26382, 26021, 25414, 
    24706, 23936,
  26863, 26824, 26760, 26638, 26065, 25008, 23662, 22893, 22516, 22526, 
    22752, 23399, 24320, 25625, 26631, 26997, 26823, 26375, 26021, 25495, 
    24769, 24164,
  26644, 26591, 26679, 26579, 26073, 25053, 23658, 22943, 22536, 22572, 
    22846, 23370, 24174, 25518, 26713, 26991, 26948, 26482, 26063, 25569, 
    24858, 24230,
  26446, 26391, 26669, 26529, 26050, 25072, 23706, 22949, 22554, 22583, 
    22942, 23426, 24396, 25301, 26357, 27031, 27029, 26510, 26110, 25612, 
    24972, 24203,
  26334, 26288, 26631, 26544, 26116, 25126, 23741, 22945, 22562, 22594, 
    22800, 23474, 24362, 25550, 26960, 27010, 26966, 26532, 26054, 25625, 
    24947, 24196,
  26319, 26292, 26588, 26565, 26107, 25083, 23762, 22993, 22606, 22643, 
    22922, 23322, 24253, 25348, 26565, 27023, 26991, 26446, 26124, 25654, 
    25035, 24403,
  26363, 26350, 26687, 26587, 26110, 25120, 23775, 23031, 22596, 22545, 
    22836, 23423, 24174, 25192, 26365, 26972, 27134, 26560, 26214, 25710, 
    25004, 24457,
  26402, 26382, 26672, 26616, 26132, 25145, 23852, 23028, 22632, 22599, 
    22842, 23438, 24233, 25301, 26446, 26934, 26922, 26431, 26131, 25679, 
    25073, 24410,
  26387, 26337, 26626, 26584, 26154, 25131, 23793, 23086, 22649, 22614, 
    22799, 23304, 24235, 25471, 26591, 26895, 26792, 26366, 26034, 25604, 
    25003, 24423,
  26307, 26220, 26600, 26543, 26084, 25167, 23883, 23062, 22657, 22656, 
    22856, 23336, 24269, 25233, 26307, 26937, 27221, 26590, 26137, 25735, 
    25175, 24671,
  26183, 26074, 26499, 26543, 26087, 25142, 23817, 23116, 22637, 22645, 
    22855, 23397, 24239, 25533, 26472, 26864, 27234, 26568, 26185, 25785, 
    25251, 24758,
  26056, 25951, 26309, 26400, 26064, 25167, 23858, 23086, 22687, 22667, 
    22827, 23371, 24207, 25191, 26526, 26722, 27121, 26532, 26241, 25779, 
    25321, 24865,
  25982, 25903, 26222, 26335, 26057, 25172, 23865, 23150, 22736, 22636, 
    22921, 23376, 24143, 25207, 26910, 26603, 27028, 26525, 26151, 25766, 
    25365, 24945,
  26026, 25982, 26310, 26368, 26041, 25152, 23913, 23133, 22698, 22658, 
    22841, 23374, 24148, 25070, 26550, 26650, 26891, 26351, 26068, 25722, 
    25308, 25072,
  26230, 26214, 26526, 26494, 26051, 25141, 23882, 23112, 22695, 22624, 
    22841, 23343, 24199, 25193, 26481, 26734, 26822, 26307, 25992, 25635, 
    25346, 24925,
  26562, 26559, 26823, 26610, 26135, 25175, 23879, 23109, 22712, 22630, 
    22857, 23310, 24248, 25196, 26389, 26937, 26903, 26264, 25950, 25536, 
    25117, 24898,
  26925, 26928, 26970, 26745, 26170, 25189, 23913, 23126, 22738, 22595, 
    22792, 23350, 24246, 25084, 26338, 27046, 26878, 26264, 25860, 25523, 
    25072, 24743,
  27208, 27231, 26996, 26779, 26221, 25163, 23934, 23176, 22762, 22609, 
    22892, 23347, 24058, 25130, 26485, 27065, 26859, 26192, 25784, 25405, 
    24919, 24502,
  27362, 27428, 27046, 26785, 26241, 25197, 23948, 23155, 22747, 22655, 
    22997, 23367, 24145, 25074, 26673, 27026, 26454, 26018, 25735, 25298, 
    24893, 24488,
  27408, 27520, 27060, 26782, 26212, 25219, 23934, 23197, 22694, 22692, 
    22954, 23256, 24216, 25260, 26143, 27001, 26685, 26082, 25673, 25255, 
    24816, 24528,
  27393, 27519, 27059, 26774, 26238, 25228, 23958, 23176, 22759, 22701, 
    22914, 23408, 24127, 25621, 26532, 27043, 26822, 26170, 25735, 25255, 
    24803, 24495,
  27329, 27424, 27014, 26742, 26235, 25194, 23954, 23217, 22782, 22606, 
    22843, 23395, 24147, 25293, 26316, 26968, 26703, 26134, 25694, 25330, 
    24816, 24421,
  27180, 27220, 27079, 26774, 26264, 25239, 23968, 23217, 22784, 22634, 
    22922, 23370, 24283, 25365, 26595, 26963, 26572, 25903, 25604, 25161, 
    24701, 24387,
  26896, 26888, 26957, 26782, 26278, 25211, 23958, 23232, 22817, 22671, 
    22840, 23415, 24196, 25353, 26367, 26943, 26965, 26148, 25701, 25199, 
    24708, 24206,
  26460, 26428, 26782, 26675, 26232, 25233, 24020, 23217, 22773, 22700, 
    22925, 23349, 24277, 25388, 26420, 26915, 26678, 25910, 25507, 25055, 
    24567, 24226,
  25898, 25871, 26506, 26516, 26154, 25289, 23930, 23173, 22826, 22703, 
    22859, 23357, 24285, 25376, 26250, 26595, 26473, 25866, 25507, 25105, 
    24637, 24179,
  25271, 25269, 26084, 26276, 26046, 25247, 23971, 23252, 22799, 22746, 
    22933, 23387, 24156, 25286, 26464, 26191, 26622, 26082, 25659, 25149, 
    24618, 24105,
  24669, 24698, 25793, 26054, 25969, 25216, 23992, 23228, 22831, 22657, 
    22913, 23380, 24119, 25211, 26260, 25854, 26603, 26235, 25776, 25223, 
    24784, 24266,
  24201, 24250, 25600, 25925, 25928, 25174, 24003, 23225, 22831, 22717, 
    22808, 23344, 23996, 25348, 26575, 25548, 26672, 26422, 25970, 25372, 
    24854, 24367,
  23949, 23997, 25453, 25907, 25960, 25211, 23975, 23249, 22813, 22692, 
    22896, 23380, 24262, 25381, 26435, 25389, 26660, 26690, 26164, 25547, 
    24867, 24306,
  23922, 23953, 25613, 25995, 25966, 25211, 23992, 23220, 22790, 22743, 
    22916, 23334, 24159, 25418, 26571, 25582, 26903, 26762, 26343, 25659, 
    24994, 24494,
  24038, 24061, 25887, 26157, 26007, 25233, 23985, 23217, 22863, 22714, 
    22942, 23354, 24218, 25178, 26223, 25988, 27226, 26784, 26247, 25703, 
    25071, 24534,
  24166, 24208, 26079, 26206, 26026, 25264, 23947, 23235, 22881, 22712, 
    22928, 23385, 24149, 25218, 26619, 26204, 27345, 26813, 26329, 25776, 
    25007, 24494,
  24192, 24263, 26034, 26241, 26049, 25219, 23965, 23235, 22831, 22749, 
    22962, 23435, 24297, 25341, 26262, 26317, 27276, 26899, 26295, 25671, 
    24962, 24434,
  24056, 24140, 25976, 26151, 26007, 25227, 23937, 23211, 22781, 22758, 
    22899, 23301, 24295, 25362, 26539, 26267, 27207, 26842, 26295, 25726, 
    25045, 24534,
  23753, 23835, 25854, 26128, 25937, 25174, 23947, 23211, 22866, 22706, 
    22957, 23199, 24262, 25218, 26579, 26242, 27276, 26820, 26316, 25796, 
    25020, 24534,
  23311, 23409, 25463, 25823, 25814, 25115, 23923, 23193, 22831, 22752, 
    22931, 23385, 24127, 25248, 26714, 25882, 27289, 26892, 26350, 25796, 
    25084, 24554,
  22783, 22924, 24926, 25484, 25668, 25093, 23930, 23211, 22861, 22735, 
    22897, 23385, 24231, 25367, 26826, 25206, 26685, 26726, 26316, 25771, 
    25090, 24501,
  22236, 22420, 24570, 25176, 25502, 25012, 23899, 23229, 22866, 22778, 
    22945, 23398, 24127, 25339, 26579, 24729, 26354, 26596, 26260, 25740, 
    25154, 24454,
  21735, 21942, 24231, 25001, 25399, 24958, 23902, 23214, 22843, 22784, 
    22982, 23342, 24164, 25244, 26537, 24300, 25999, 26539, 26232, 25684, 
    25014, 24401,
  21347, 21557, 23969, 24818, 25313, 24922, 23882, 23247, 22899, 22752, 
    22871, 23357, 24219, 25421, 26406, 23821, 25956, 26582, 26247, 25834, 
    25097, 24582,
  21130, 21330, 23858, 24778, 25285, 24894, 23889, 23203, 22858, 22819, 
    22985, 23459, 24201, 25188, 26573, 23640, 25850, 26610, 26301, 25853, 
    25186, 24669,
  21119, 21300, 24051, 24843, 25293, 24869, 23850, 23197, 22881, 22767, 
    23051, 23413, 24290, 25167, 26504, 23849, 25881, 26597, 26316, 25926, 
    25224, 24649,
  21302, 21471, 24221, 24934, 25331, 24920, 23865, 23161, 22870, 22813, 
    22966, 23467, 24374, 25153, 26549, 24141, 26043, 26597, 26329, 25971, 
    25206, 24669,
  21619, 21795, 24208, 24953, 25351, 24908, 23802, 23183, 22867, 22787, 
    22940, 23340, 24256, 25316, 26507, 24107, 25906, 26503, 26301, 25840, 
    25161, 24670,
  21993, 22165, 24190, 24999, 25339, 24880, 23820, 23203, 22900, 22879, 
    22926, 23379, 24271, 25272, 26822, 23993, 25800, 26568, 26323, 25903, 
    25276, 24730,
  22340, 22475, 24518, 25145, 25393, 24900, 23837, 23171, 22888, 22834, 
    23032, 23422, 24234, 25300, 26350, 24213, 25888, 26560, 26329, 25891, 
    25270, 24764,
  22588, 22679, 24675, 25255, 25425, 24867, 23820, 23206, 22897, 22820, 
    22975, 23353, 24286, 25403, 26591, 24346, 25943, 26496, 26248, 25791, 
    25200, 24697,
  22700, 22785, 24723, 25242, 25403, 24794, 23792, 23189, 22882, 22805, 
    23024, 23536, 24296, 25089, 26532, 24348, 25881, 26525, 26206, 25841, 
    25168, 24670,
  22686, 22793, 24584, 25161, 25388, 24833, 23757, 23175, 22880, 22837, 
    22998, 23529, 24333, 25342, 26795, 24296, 26018, 26503, 26193, 25667, 
    25143, 24637,
  22558, 22671, 24503, 25177, 25377, 24760, 23734, 23157, 22895, 22892, 
    23069, 23473, 24235, 25368, 26532, 24326, 26018, 26453, 26226, 25704, 
    25201, 24731,
  22299, 22389, 24577, 25153, 25322, 24769, 23734, 23160, 22883, 22938, 
    22941, 23478, 24309, 25347, 26882, 24470, 26087, 26496, 26207, 25748, 
    25258, 24738,
  21895, 21969, 24318, 25019, 25294, 24758, 23765, 23157, 22907, 22915, 
    23036, 23550, 24410, 25417, 26535, 24289, 26044, 26518, 26110, 25704, 
    25207, 24738,
  21411, 21511, 24064, 24817, 25185, 24716, 23734, 23149, 22904, 22904, 
    23064, 23474, 24235, 25517, 26601, 23968, 25907, 26460, 26117, 25624, 
    25131, 24651,
  21009, 21163, 23852, 24723, 25220, 24702, 23724, 23155, 22919, 22881, 
    23022, 23568, 24302, 25461, 26689, 23753, 25751, 26403, 26014, 25531, 
    25080, 24585,
  20866, 21058, 23819, 24693, 25117, 24685, 23696, 23143, 22925, 22973, 
    23096, 23538, 24401, 25454, 26956, 23756, 25857, 26317, 25897, 25482, 
    24972, 24431,
  21039, 21232, 23934, 24718, 25117, 24646, 23640, 23152, 22911, 22907, 
    23014, 23525, 24465, 25346, 26468, 23931, 25914, 26288, 25951, 25506, 
    24858, 24471,
  21428, 21605, 24144, 24853, 25174, 24615, 23644, 23123, 22914, 22899, 
    23034, 23589, 24418, 25406, 26881, 24190, 25976, 26338, 26014, 25519, 
    24966, 24605,
  21846, 22029, 24344, 24995, 25175, 24613, 23603, 23126, 22873, 22988, 
    23063, 23584, 24320, 25404, 26713, 24398, 25976, 26317, 26056, 25644, 
    25043, 24512,
  22143, 22356, 24535, 25117, 25183, 24605, 23596, 23097, 22961, 22986, 
    23162, 23656, 24362, 25607, 26829, 24590, 25989, 26281, 26015, 25520, 
    24954, 24492,
  22275, 22511, 24659, 25144, 25226, 24569, 23607, 23121, 22929, 22908, 
    23120, 23653, 24481, 25558, 26813, 24676, 26095, 26296, 26029, 25495, 
    24853, 24519,
  22292, 22527, 24662, 25111, 25212, 24535, 23607, 23085, 22959, 22929, 
    23126, 23595, 24375, 25653, 26626, 24553, 26064, 26353, 26091, 25564, 
    25044, 24479,
  22285, 22502, 24629, 25128, 25207, 24516, 23558, 23127, 22944, 22898, 
    23092, 23679, 24301, 25616, 26920, 24419, 25907, 26339, 26057, 25620, 
    25108, 24654,
  22311, 22506, 24639, 25141, 25161, 24505, 23524, 23083, 22944, 23035, 
    23058, 23763, 24452, 25465, 26816, 24380, 25907, 26354, 26084, 25726, 
    25191, 24547,
  22375, 22541, 24652, 25196, 25167, 24424, 23531, 23086, 22947, 23021, 
    23121, 23621, 24506, 25819, 26826, 24355, 25951, 26289, 26071, 25714, 
    25095, 24627,
  22457, 22588, 24688, 25166, 25124, 24373, 23476, 23078, 22977, 23033, 
    23141, 23700, 24452, 25647, 26743, 24290, 25959, 26282, 26078, 25565, 
    25115, 24588,
  22554, 22653, 24772, 25193, 25139, 24373, 23455, 23072, 22942, 22967, 
    23139, 23673, 24534, 25901, 26889, 24323, 25965, 26268, 26037, 25626, 
    25007, 24575,
  22690, 22764, 24871, 25228, 25119, 24320, 23459, 23075, 23021, 23005, 
    23153, 23701, 24534, 25798, 26671, 24442, 26034, 26254, 25920, 25540, 
    24905, 24300,
  22896, 22946, 25023, 25325, 25079, 24304, 23442, 23105, 22975, 22985, 
    23171, 23815, 24478, 25737, 26945, 24576, 26270, 26225, 25969, 25584, 
    24989, 24408,
  23183, 23206, 25155, 25368, 25054, 24259, 23376, 23067, 22981, 23085, 
    23151, 23686, 24552, 25954, 26913, 24740, 26226, 26247, 25948, 25578, 
    24932, 24489,
  23516, 23517, 25238, 25409, 25028, 24175, 23384, 23088, 22967, 23054, 
    23052, 23742, 24582, 25607, 26860, 24829, 26171, 26153, 25914, 25454, 
    24913, 24435,
  23842, 23823, 25365, 25369, 25025, 24156, 23332, 23050, 23046, 22983, 
    23200, 23702, 24737, 25976, 26875, 24809, 26140, 26168, 25804, 25355, 
    24780, 24248,
  24139, 24086, 25333, 25471, 24980, 24103, 23328, 23071, 22985, 22989, 
    23152, 23674, 24530, 25906, 26715, 24535, 26022, 26082, 25763, 25355, 
    24741, 24262,
  24386, 24286, 25356, 25348, 24931, 24047, 23339, 23065, 23032, 23041, 
    23198, 23814, 24637, 26029, 26860, 24359, 25823, 26032, 25728, 25269, 
    24742, 24289,
  24494, 24356, 25275, 25342, 24834, 23994, 23256, 23018, 23044, 23030, 
    23249, 23763, 24851, 26019, 27204, 24320, 25848, 25996, 25619, 25175, 
    24729, 24182,
  24368, 24221, 25331, 25299, 24800, 23941, 23242, 23086, 22986, 23102, 
    23281, 23857, 24768, 26222, 27047, 24344, 25873, 25895, 25550, 25095, 
    24602, 24122,
  24096, 23960, 25320, 25251, 24729, 23905, 23221, 23034, 23039, 23025, 
    23324, 23837, 24952, 26289, 27057, 24433, 25848, 25845, 25522, 25089, 
    24431, 24116,
  23953, 23824, 25354, 25294, 24652, 23799, 23187, 23037, 23009, 23111, 
    23298, 23850, 24933, 26282, 27174, 24567, 26029, 25773, 25399, 24916, 
    24406, 23889,
  27893, 27823, 27182, 26597, 25522, 24109, 22734, 22246, 22179, 22498, 
    22895, 23699, 24612, 25893, 26806, 27575, 26866, 25929, 25433, 24831, 
    24216, 23758,
  27840, 27770, 27132, 26670, 25576, 24190, 22803, 22308, 22167, 22580, 
    22943, 23661, 24593, 25635, 26466, 27576, 27015, 26046, 25537, 25024, 
    24305, 23704,
  27731, 27666, 26894, 26484, 25596, 24274, 22910, 22319, 22158, 22514, 
    22866, 23508, 24496, 25685, 26543, 27259, 26878, 26117, 25564, 25049, 
    24228, 23804,
  27648, 27597, 26787, 26435, 25584, 24332, 22972, 22360, 22216, 22540, 
    22845, 23579, 24457, 25751, 26597, 26840, 26324, 25843, 25474, 25005, 
    24247, 23744,
  27622, 27579, 26724, 26368, 25598, 24388, 23049, 22484, 22230, 22513, 
    22973, 23518, 24503, 25848, 26592, 26676, 25839, 25620, 25336, 24849, 
    24183, 23569,
  27623, 27569, 26949, 26513, 25676, 24464, 23107, 22481, 22263, 22585, 
    22822, 23536, 24537, 25779, 26403, 26866, 26423, 25785, 25377, 24780, 
    24157, 23602,
  27614, 27550, 27106, 26710, 25888, 24528, 23177, 22513, 22333, 22533, 
    22936, 23457, 24510, 25816, 26822, 27251, 26890, 25929, 25342, 24755, 
    24176, 23716,
  27579, 27536, 27207, 26849, 25956, 24620, 23214, 22568, 22311, 22530, 
    22844, 23538, 24530, 25520, 26684, 27469, 27051, 25885, 25349, 24811, 
    24169, 23682,
  27520, 27519, 27201, 26839, 26001, 24659, 23239, 22571, 22311, 22544, 
    22907, 23525, 24384, 25629, 26625, 27553, 26747, 25749, 25259, 24760, 
    24137, 23662,
  27444, 27467, 27179, 26860, 26053, 24751, 23325, 22636, 22367, 22538, 
    22892, 23499, 24480, 25790, 26969, 27567, 26709, 25726, 25231, 24630, 
    24067, 23655,
  27345, 27371, 27182, 26829, 26047, 24751, 23352, 22632, 22366, 22552, 
    22863, 23511, 24467, 25715, 26598, 27503, 26821, 25942, 25417, 24773, 
    24162, 23681,
  27217, 27259, 27142, 26798, 26050, 24804, 23435, 22673, 22389, 22543, 
    22835, 23595, 24479, 25566, 26744, 27420, 26907, 26129, 25575, 24978, 
    24174, 23694,
  27080, 27153, 27081, 26739, 26026, 24844, 23449, 22753, 22386, 22525, 
    22780, 23313, 24354, 25601, 26282, 27378, 26982, 26332, 25809, 25114, 
    24345, 23834,
  26983, 27063, 26944, 26696, 26006, 24877, 23494, 22758, 22430, 22514, 
    22777, 23521, 24351, 25613, 26423, 27356, 27188, 26476, 25932, 25294, 
    24435, 23860,
  26958, 27004, 26875, 26657, 26047, 24955, 23532, 22773, 22424, 22508, 
    22908, 23495, 24284, 25510, 26659, 27359, 27194, 26510, 26064, 25412, 
    24581, 23961,
  26992, 26991, 26938, 26695, 26066, 24938, 23553, 22837, 22450, 22568, 
    22873, 23497, 24244, 25177, 26249, 27307, 27126, 26540, 26037, 25393, 
    24568, 23927,
  27043, 27015, 27029, 26671, 26101, 25000, 23587, 22849, 22473, 22553, 
    22881, 23411, 24353, 25452, 26551, 27284, 27069, 26417, 25974, 25337, 
    24586, 23960,
  27067, 27023, 26981, 26668, 26129, 25000, 23629, 22919, 22511, 22613, 
    22836, 23456, 24330, 25261, 26348, 27242, 27113, 26554, 26174, 25486, 
    24643, 24027,
  27025, 26961, 26901, 26690, 26095, 25041, 23646, 22907, 22534, 22601, 
    22884, 23418, 24246, 25463, 26735, 27228, 27088, 26604, 26201, 25672, 
    24860, 24214,
  26901, 26822, 26844, 26646, 26076, 25033, 23660, 22901, 22545, 22621, 
    22904, 23402, 24268, 25449, 26821, 27091, 26976, 26554, 26125, 25715, 
    24917, 24274,
  26727, 26658, 26806, 26603, 26149, 25021, 23722, 22919, 22539, 22580, 
    22932, 23341, 24150, 25502, 26575, 27089, 26932, 26575, 26229, 25740, 
    25069, 24414,
  26574, 26539, 26788, 26609, 26091, 25091, 23770, 22954, 22603, 22552, 
    22929, 23382, 24201, 25398, 26328, 27075, 26963, 26604, 26256, 25759, 
    25050, 24367,
  26504, 26504, 26679, 26603, 26085, 25108, 23718, 23021, 22612, 22594, 
    22815, 23402, 24208, 25393, 26548, 27085, 27069, 26590, 26194, 25746, 
    25024, 24380,
  26527, 26539, 26682, 26609, 26126, 25142, 23773, 23009, 22623, 22609, 
    22897, 23452, 24117, 25504, 26707, 27031, 27225, 26647, 26214, 25751, 
    25094, 24380,
  26596, 26596, 26807, 26641, 26128, 25097, 23763, 23036, 22597, 22617, 
    22914, 23452, 24215, 25414, 26522, 27035, 26963, 26510, 26221, 25757, 
    25049, 24541,
  26644, 26620, 26884, 26665, 26140, 25130, 23832, 23044, 22632, 22640, 
    22854, 23305, 24343, 25325, 26864, 27120, 27038, 26546, 26097, 25626, 
    25011, 24507,
  26617, 26574, 26740, 26635, 26114, 25099, 23846, 23071, 22746, 22700, 
    22908, 23411, 24195, 25313, 26482, 27092, 27181, 26501, 26138, 25664, 
    25074, 24594,
  26507, 26456, 26710, 26576, 26140, 25150, 23839, 23091, 22666, 22642, 
    22868, 23497, 24195, 25364, 26451, 26970, 27144, 26574, 26138, 25720, 
    25080, 24674,
  26336, 26285, 26559, 26519, 26091, 25130, 23811, 23112, 22725, 22636, 
    22853, 23375, 24281, 25360, 26689, 26875, 27037, 26459, 26138, 25720, 
    25208, 24848,
  26142, 26101, 26422, 26414, 26107, 25119, 23904, 23126, 22716, 22667, 
    22936, 23415, 24215, 25443, 26235, 26700, 27031, 26466, 26138, 25757, 
    25278, 24935,
  25981, 25962, 26331, 26385, 26042, 25174, 23880, 23143, 22727, 22641, 
    22859, 23369, 24165, 25534, 26839, 26654, 26838, 26372, 26075, 25701, 
    25341, 24955,
  25932, 25934, 26354, 26363, 26071, 25110, 23866, 23132, 22727, 22699, 
    22856, 23415, 24231, 25357, 26506, 26657, 26888, 26271, 25999, 25645, 
    25277, 24935,
  26062, 26066, 26384, 26384, 26042, 25132, 23935, 23164, 22759, 22601, 
    22867, 23364, 24369, 25227, 26409, 26685, 26938, 26285, 25923, 25545, 
    25073, 24821,
  26367, 26351, 26682, 26635, 26171, 25174, 23904, 23176, 22768, 22698, 
    22881, 23389, 24258, 25457, 26388, 26865, 26919, 26242, 25826, 25483, 
    24952, 24660,
  26757, 26725, 27018, 26788, 26204, 25197, 23921, 23158, 22756, 22626, 
    22898, 23557, 24093, 25224, 26659, 27110, 26912, 26213, 25826, 25358, 
    24830, 24478,
  27114, 27092, 27069, 26826, 26271, 25267, 23949, 23187, 22729, 22692, 
    22880, 23402, 24181, 25494, 26599, 27151, 26918, 26226, 25785, 25389, 
    24786, 24505,
  27357, 27371, 27089, 26753, 26254, 25233, 23897, 23151, 22779, 22701, 
    22961, 23381, 24226, 25361, 26301, 27124, 26719, 26097, 25778, 25345, 
    24849, 24411,
  27463, 27519, 27122, 26807, 26257, 25255, 23921, 23154, 22811, 22617, 
    22997, 23391, 24092, 25350, 26785, 27110, 26956, 26226, 25798, 25382, 
    24753, 24377,
  27444, 27520, 27072, 26823, 26291, 25258, 23962, 23222, 22776, 22720, 
    22900, 23404, 24282, 25559, 26632, 27207, 27081, 26292, 25826, 25376, 
    24811, 24364,
  27300, 27361, 27109, 26896, 26262, 25272, 23935, 23184, 22855, 22712, 
    22920, 23416, 24124, 25280, 26249, 27207, 27179, 26335, 25895, 25339, 
    24906, 24431,
  27002, 27021, 27101, 26882, 26317, 25297, 23966, 23181, 22785, 22648, 
    22954, 23386, 24221, 25280, 26297, 27126, 27062, 26270, 25757, 25283, 
    24677, 24303,
  26517, 26493, 26840, 26794, 26234, 25241, 23952, 23255, 22817, 22726, 
    22900, 23431, 24176, 25194, 26538, 26987, 26781, 26110, 25625, 25133, 
    24658, 24263,
  25858, 25809, 26549, 26578, 26196, 25264, 23969, 23166, 22811, 22737, 
    22886, 23394, 24205, 25405, 26521, 26698, 26625, 25872, 25501, 25139, 
    24645, 24269,
  25099, 25050, 26101, 26222, 26026, 25210, 23955, 23234, 22846, 22692, 
    22983, 23467, 24035, 25324, 26476, 26107, 26538, 26032, 25632, 25220, 
    24638, 24256,
  24356, 24326, 25577, 25893, 25938, 25202, 23955, 23207, 22796, 22740, 
    22882, 23373, 24119, 25338, 26169, 25542, 26538, 26465, 25929, 25326, 
    24753, 24437,
  23746, 23743, 25412, 25821, 25910, 25171, 23972, 23201, 22872, 22783, 
    22925, 23406, 24228, 25259, 26521, 25286, 26625, 26718, 26232, 25494, 
    24906, 24363,
  23358, 23380, 25239, 25672, 25847, 25165, 23959, 23204, 22843, 22737, 
    23005, 23409, 24190, 25163, 26365, 25150, 26725, 26819, 26274, 25643, 
    24995, 24451,
  23222, 23250, 25115, 25624, 25824, 25151, 23945, 23207, 22820, 22723, 
    22957, 23347, 24149, 25321, 26382, 24980, 26837, 26848, 26406, 25712, 
    24951, 24484,
  23286, 23293, 25062, 25599, 25806, 25157, 23965, 23219, 22828, 22737, 
    22954, 23363, 24205, 25333, 26454, 25019, 26837, 26841, 26371, 25860, 
    25072, 24591,
  23416, 23398, 25166, 25707, 25784, 25145, 23997, 23227, 22840, 22755, 
    23011, 23360, 24104, 25417, 26367, 25164, 26956, 26870, 26364, 25779, 
    25021, 24544,
  23456, 23442, 25252, 25667, 25784, 25134, 23952, 23234, 22826, 22752, 
    22954, 23353, 24269, 25212, 26251, 25283, 26781, 26782, 26343, 25718, 
    25033, 24464,
  23316, 23330, 25176, 25604, 25751, 25106, 23938, 23181, 22878, 22766, 
    23028, 23327, 24129, 25354, 26257, 25172, 26825, 26826, 26357, 25724, 
    25002, 24397,
  22996, 23035, 24902, 25457, 25643, 25103, 23917, 23195, 22902, 22743, 
    22891, 23358, 24119, 25159, 26593, 24913, 26526, 26768, 26378, 25712, 
    24976, 24457,
  22557, 22611, 24570, 25212, 25544, 25084, 23966, 23204, 22840, 22775, 
    22991, 23482, 24267, 25249, 26513, 24632, 26239, 26703, 26323, 25768, 
    25008, 24471,
  22074, 22153, 24197, 24972, 25437, 24994, 23893, 23260, 22834, 22763, 
    22909, 23384, 24144, 25324, 26523, 24234, 26007, 26653, 26254, 25743, 
    25015, 24498,
  21623, 21742, 24020, 24843, 25346, 25003, 23952, 23255, 22864, 22829, 
    23057, 23439, 24282, 25475, 26775, 23841, 25840, 26573, 26316, 25799, 
    25002, 24444,
  21272, 21424, 23900, 24829, 25317, 24944, 23876, 23181, 22852, 22801, 
    23026, 23523, 24250, 25303, 26610, 23844, 25982, 26566, 26323, 25787, 
    25085, 24464,
  21067, 21228, 23837, 24770, 25329, 24941, 23903, 23237, 22870, 22781, 
    22966, 23490, 24134, 25345, 26632, 23771, 25921, 26610, 26385, 25799, 
    25244, 24599,
  21019, 21177, 23890, 24773, 25317, 24930, 23903, 23228, 22896, 22812, 
    23006, 23450, 24112, 25370, 26594, 23682, 25790, 26682, 26385, 25935, 
    25251, 24679,
  21116, 21265, 24126, 24864, 25338, 24896, 23872, 23181, 22914, 22850, 
    22989, 23389, 24132, 25341, 26470, 23857, 25865, 26675, 26413, 25912, 
    25238, 24800,
  21331, 21468, 24276, 24986, 25326, 24871, 23848, 23205, 22885, 22790, 
    22969, 23511, 24211, 25403, 26103, 24085, 26065, 26632, 26441, 25900, 
    25283, 24760,
  21624, 21756, 24385, 25002, 25372, 24913, 23844, 23173, 22902, 22816, 
    22943, 23493, 24322, 25450, 26594, 24182, 26046, 26610, 26413, 25912, 
    25271, 24713,
  21948, 22086, 24292, 24978, 25398, 24911, 23866, 23211, 22873, 22822, 
    22992, 23351, 24327, 25548, 26540, 24043, 25791, 26567, 26337, 25918, 
    25220, 24680,
  22263, 22398, 24436, 25042, 25355, 24835, 23817, 23179, 22897, 22833, 
    23030, 23478, 24394, 25397, 26524, 24098, 25822, 26531, 26365, 25812, 
    25239, 24666,
  22539, 22640, 24576, 25134, 25410, 24880, 23786, 23167, 22885, 22879, 
    23061, 23514, 24322, 25166, 26285, 24218, 25847, 26545, 26303, 25850, 
    25245, 24754,
  22742, 22803, 24644, 25159, 25430, 24849, 23755, 23149, 22859, 22859, 
    23044, 23476, 24224, 25301, 26492, 24282, 25853, 26574, 26345, 25844, 
    25252, 24788,
  22838, 22893, 24695, 25180, 25396, 24838, 23776, 23155, 22900, 22848, 
    23107, 23405, 24303, 25364, 26315, 24296, 25897, 26560, 26282, 25794, 
    25265, 24834,
  22806, 22888, 24596, 25175, 25381, 24782, 23769, 23165, 22901, 22805, 
    23116, 23515, 24308, 25648, 26438, 24370, 25990, 26589, 26200, 25820, 
    25176, 24754,
  22636, 22733, 24657, 25153, 25355, 24802, 23755, 23186, 22901, 22880, 
    23021, 23487, 24276, 25467, 26720, 24515, 26072, 26517, 26179, 25707, 
    25189, 24708,
  22314, 22397, 24701, 25224, 25347, 24721, 23728, 23150, 22924, 22909, 
    23033, 23561, 24276, 25518, 26665, 24629, 26209, 26481, 26193, 25764, 
    25176, 24788,
  21855, 21926, 24564, 25100, 25290, 24732, 23714, 23142, 22930, 22932, 
    23070, 23500, 24353, 25488, 26701, 24486, 26084, 26445, 26131, 25632, 
    25081, 24601,
  21350, 21453, 24194, 24976, 25270, 24710, 23728, 23177, 22916, 22898, 
    23059, 23482, 24173, 25365, 26706, 24149, 25979, 26387, 26097, 25701, 
    25030, 24581,
  20973, 21149, 23963, 24796, 25190, 24696, 23662, 23142, 22907, 22930, 
    23068, 23465, 24346, 25509, 26539, 23979, 25935, 26401, 26014, 25503, 
    24935, 24554,
  20886, 21120, 23928, 24721, 25141, 24654, 23683, 23160, 22902, 22967, 
    23088, 23450, 24484, 25553, 26517, 23858, 25904, 26316, 26007, 25485, 
    24935, 24441,
  21119, 21356, 23938, 24818, 25156, 24635, 23670, 23163, 22905, 22896, 
    23043, 23529, 24369, 25601, 26898, 23936, 25823, 26309, 26063, 25628, 
    25024, 24575,
  21554, 21756, 24237, 24963, 25193, 24626, 23638, 23110, 22925, 22933, 
    23077, 23491, 24371, 25660, 26785, 24189, 25942, 26395, 26056, 25597, 
    24987, 24535,
  22006, 22185, 24483, 25044, 25242, 24593, 23635, 23140, 22949, 22896, 
    23063, 23572, 24394, 25514, 26804, 24421, 25935, 26359, 26035, 25628, 
    25012, 24509,
  22333, 22521, 24649, 25141, 25222, 24604, 23597, 23152, 22955, 23002, 
    23027, 23586, 24487, 25704, 27056, 24615, 26023, 26351, 26029, 25610, 
    24981, 24429,
  22487, 22690, 24681, 25128, 25214, 24574, 23594, 23111, 22941, 22986, 
    23141, 23614, 24387, 25577, 26889, 24682, 26167, 26367, 26071, 25629, 
    25019, 24509,
  22507, 22711, 24570, 25128, 25162, 24478, 23598, 23117, 22947, 22934, 
    23115, 23560, 24444, 25768, 26850, 24489, 25960, 26338, 26084, 25747, 
    24988, 24610,
  22482, 22673, 24581, 25112, 25197, 24493, 23518, 23144, 22953, 22989, 
    23141, 23596, 24461, 25589, 26954, 24332, 25793, 26353, 26106, 25754, 
    25128, 24644,
  22476, 22650, 24667, 25118, 25191, 24448, 23511, 23091, 22939, 23064, 
    23210, 23673, 24550, 25798, 26887, 24360, 25849, 26339, 26106, 25710, 
    25065, 24644,
  22499, 22653, 24730, 25199, 25217, 24434, 23497, 23088, 22954, 23041, 
    23139, 23592, 24499, 25668, 27025, 24446, 26017, 26310, 26078, 25654, 
    25148, 24644,
  22530, 22668, 24789, 25166, 25117, 24429, 23480, 23112, 22948, 22981, 
    23191, 23668, 24600, 25548, 26651, 24432, 25949, 26353, 26113, 25673, 
    25072, 24578,
  22573, 22702, 24847, 25226, 25077, 24347, 23418, 23086, 22975, 22976, 
    23125, 23666, 24612, 25769, 26882, 24467, 26043, 26303, 25975, 25593, 
    25059, 24471,
  22663, 22787, 24913, 25242, 25097, 24295, 23467, 23086, 22960, 23053, 
    23142, 23646, 24561, 25673, 26846, 24674, 26199, 26289, 25920, 25544, 
    24926, 24397,
  22847, 22955, 24982, 25323, 25080, 24219, 23384, 23075, 22993, 23040, 
    23146, 23669, 24583, 25934, 26766, 24771, 26204, 26310, 25941, 25599, 
    25028, 24525,
  23137, 23218, 25179, 25337, 25072, 24228, 23391, 23102, 22973, 22991, 
    23203, 23687, 24593, 25781, 26734, 24798, 26199, 26253, 25914, 25463, 
    24920, 24432,
  23494, 23546, 25253, 25407, 25040, 24183, 23367, 23099, 23019, 23000, 
    23146, 23705, 24660, 25843, 26928, 24873, 26168, 26167, 25825, 25470, 
    24831, 24418,
  23849, 23870, 25380, 25450, 24992, 24136, 23343, 23090, 23026, 22997, 
    23218, 23779, 24835, 26126, 27067, 24848, 26124, 26131, 25832, 25364, 
    24774, 24318,
  24159, 24137, 25408, 25404, 24972, 24156, 23360, 23082, 23035, 23124, 
    23255, 23720, 24715, 26113, 27129, 24540, 25907, 26117, 25776, 25296, 
    24825, 24366,
  24398, 24319, 25319, 25351, 24892, 24122, 23319, 23070, 23003, 23092, 
    23253, 23838, 24782, 26123, 26499, 24217, 25726, 26088, 25776, 25402, 
    24775, 24453,
  24494, 24366, 25322, 25318, 24855, 24030, 23260, 23109, 23076, 23116, 
    23273, 23795, 24915, 26114, 27465, 24091, 25764, 25979, 25639, 25247, 
    24839, 24306,
  24371, 24223, 25328, 25262, 24779, 24002, 23303, 23088, 23056, 23093, 
    23281, 23904, 24787, 26092, 26946, 23967, 25565, 25887, 25584, 25166, 
    24636, 24253,
  24116, 23972, 25239, 25257, 24716, 23856, 23268, 23095, 23068, 23102, 
    23301, 23869, 24920, 26210, 27419, 24053, 25584, 25851, 25537, 25160, 
    24616, 24153,
  23983, 23844, 25302, 25257, 24664, 23871, 23202, 23101, 23048, 23079, 
    23322, 23971, 24918, 26181, 27307, 24299, 25851, 25743, 25489, 25049, 
    24477, 23952,
  27903, 27799, 27198, 26574, 25518, 24057, 22739, 22289, 22175, 22558, 
    22930, 23616, 24641, 25728, 26887, 27601, 26841, 26010, 25429, 24912, 
    24221, 23700,
  27850, 27754, 27120, 26625, 25604, 24161, 22833, 22303, 22140, 22558, 
    22918, 23702, 24762, 25621, 26756, 27654, 27109, 26082, 25546, 24974, 
    24335, 23653,
  27737, 27666, 26963, 26499, 25601, 24247, 22926, 22327, 22180, 22552, 
    22881, 23659, 24816, 25807, 26671, 27335, 26903, 26089, 25525, 24955, 
    24271, 23727,
  27651, 27611, 26889, 26467, 25626, 24354, 22978, 22430, 22257, 22600, 
    22872, 23623, 24599, 25891, 26707, 27065, 26492, 25923, 25477, 24918, 
    24303, 23559,
  27624, 27597, 26909, 26515, 25693, 24409, 23051, 22406, 22262, 22519, 
    22860, 23562, 24552, 25725, 26634, 27065, 26529, 25835, 25290, 24768, 
    24112, 23505,
  27628, 27587, 27087, 26646, 25787, 24535, 23144, 22500, 22300, 22548, 
    22849, 23587, 24453, 25739, 26607, 27310, 26754, 25764, 25242, 24650, 
    24041, 23464,
  27622, 27572, 27244, 26785, 25898, 24557, 23183, 22479, 22343, 22542, 
    22939, 23543, 24490, 25614, 26982, 27481, 26479, 25418, 25021, 24556, 
    24086, 23477,
  27593, 27563, 27254, 26856, 25975, 24667, 23227, 22547, 22355, 22550, 
    22942, 23589, 24541, 25818, 26571, 27557, 26423, 25468, 25000, 24556, 
    24149, 23564,
  27547, 27544, 27219, 26865, 25998, 24711, 23296, 22611, 22369, 22573, 
    22905, 23553, 24512, 25534, 26915, 27560, 26616, 25662, 25138, 24711, 
    24155, 23530,
  27485, 27481, 27182, 26891, 26078, 24725, 23359, 22596, 22357, 22538, 
    22916, 23499, 24566, 25555, 26464, 27607, 26872, 26022, 25406, 24903, 
    24142, 23731,
  27392, 27378, 27226, 26873, 26051, 24770, 23334, 22684, 22371, 22460, 
    22845, 23522, 24420, 25643, 26451, 27574, 26965, 26174, 25564, 25052, 
    24249, 23683,
  27255, 27267, 27188, 26878, 26092, 24828, 23414, 22719, 22427, 22523, 
    22810, 23481, 24385, 25555, 26389, 27519, 27026, 26310, 25757, 25127, 
    24364, 23871,
  27100, 27164, 27057, 26762, 26029, 24867, 23480, 22728, 22421, 22503, 
    22872, 23430, 24287, 25487, 26539, 27507, 27126, 26354, 25895, 25300, 
    24478, 23910,
  26979, 27064, 26976, 26707, 26009, 24909, 23469, 22760, 22406, 22609, 
    22855, 23422, 24372, 25687, 26635, 27418, 27207, 26585, 26012, 25437, 
    24631, 23963,
  26926, 26982, 26907, 26701, 26051, 24948, 23542, 22766, 22452, 22571, 
    22838, 23465, 24375, 25538, 26849, 27357, 27151, 26570, 26046, 25418, 
    24649, 23996,
  26937, 26947, 26967, 26701, 26069, 24945, 23583, 22816, 22470, 22485, 
    22923, 23404, 24281, 25600, 26444, 27307, 27151, 26504, 26039, 25467, 
    24592, 23869,
  26986, 26963, 26974, 26713, 26023, 24940, 23583, 22830, 22460, 22585, 
    22803, 23373, 24355, 25440, 26298, 27296, 27070, 26562, 26087, 25591, 
    24668, 24056,
  27036, 26987, 26951, 26685, 26054, 24973, 23663, 22895, 22551, 22596, 
    22905, 23368, 24443, 25410, 26504, 27288, 27082, 26613, 26225, 25659, 
    24846, 24237,
  27041, 26966, 26910, 26637, 26088, 25029, 23680, 22927, 22551, 22501, 
    22840, 23406, 24216, 25463, 26740, 27198, 27076, 26612, 26266, 25734, 
    25030, 24330,
  26975, 26890, 26896, 26645, 26134, 25029, 23714, 22909, 22539, 22630, 
    22842, 23390, 24393, 25133, 26468, 27140, 26895, 26554, 26210, 25765, 
    25024, 24297,
  26859, 26801, 26898, 26670, 26123, 25090, 23693, 22968, 22582, 22610, 
    22810, 23393, 24343, 25470, 26506, 27146, 27007, 26582, 26182, 25796, 
    25081, 24310,
  26757, 26752, 26826, 26679, 26079, 25079, 23752, 22982, 22602, 22569, 
    22896, 23392, 24309, 25484, 26735, 27126, 26964, 26582, 26176, 25721, 
    25081, 24256,
  26723, 26762, 26741, 26664, 26094, 25059, 23717, 22964, 22617, 22635, 
    22807, 23440, 24156, 25388, 26700, 27129, 27076, 26626, 26148, 25757, 
    25151, 24336,
  26764, 26810, 26785, 26629, 26097, 25087, 23797, 23038, 22550, 22597, 
    22821, 23425, 24218, 25520, 26298, 27104, 26988, 26575, 26210, 25776, 
    25157, 24429,
  26838, 26857, 26910, 26712, 26097, 25087, 23758, 23032, 22634, 22582, 
    22809, 23374, 24271, 25437, 26591, 27160, 26907, 26467, 26044, 25732, 
    25125, 24610,
  26884, 26870, 26879, 26685, 26128, 25109, 23800, 23087, 22660, 22585, 
    22869, 23422, 24251, 25402, 26744, 27172, 27038, 26489, 26092, 25664, 
    25169, 24596,
  26850, 26825, 26785, 26675, 26116, 25114, 23824, 23075, 22648, 22571, 
    22840, 23340, 24170, 25525, 26264, 27049, 27050, 26467, 26078, 25764, 
    25251, 24777,
  26723, 26708, 26704, 26582, 26147, 25118, 23862, 23072, 22657, 22631, 
    22806, 23436, 24365, 25357, 26503, 26868, 26764, 26423, 26147, 25745, 
    25245, 24777,
  26516, 26510, 26707, 26572, 26087, 25154, 23862, 23092, 22724, 22584, 
    22877, 23378, 24137, 25113, 26644, 26857, 26632, 26300, 26016, 25663, 
    25309, 24911,
  26252, 26251, 26778, 26542, 26110, 25151, 23886, 23089, 22768, 22647, 
    22863, 23403, 24260, 25183, 26215, 26876, 26795, 26307, 25995, 25775, 
    25264, 24884,
  25982, 25990, 26638, 26532, 26142, 25128, 23924, 23116, 22735, 22644, 
    22888, 23345, 24108, 25287, 26321, 26826, 26870, 26379, 25988, 25676, 
    25340, 24970,
  25798, 25814, 26317, 26356, 26050, 25108, 23903, 23166, 22726, 22644, 
    22799, 23413, 24085, 25178, 26775, 26634, 26863, 26373, 25954, 25613, 
    25244, 24910,
  25802, 25805, 26176, 26275, 26059, 25153, 23869, 23124, 22764, 22624, 
    22808, 23327, 24080, 25110, 26770, 26478, 26795, 26220, 25822, 25414, 
    25027, 24675,
  26029, 25999, 26438, 26445, 26119, 25190, 23899, 23192, 22770, 22641, 
    22834, 23451, 24267, 25217, 26598, 26657, 26751, 26162, 25739, 25358, 
    24893, 24461,
  26419, 26362, 26875, 26693, 26193, 25260, 23955, 23162, 22758, 22664, 
    22828, 23402, 24149, 25233, 26188, 27032, 26651, 25996, 25635, 25376, 
    24842, 24421,
  26851, 26793, 27062, 26814, 26253, 25215, 23945, 23189, 22761, 22764, 
    22913, 23456, 24124, 25450, 26556, 27159, 26676, 26082, 25704, 25264, 
    24810, 24420,
  27207, 27171, 27057, 26838, 26245, 25234, 23938, 23141, 22746, 22666, 
    22861, 23331, 24131, 25352, 26040, 27128, 26769, 26090, 25684, 25251, 
    24657, 24306,
  27406, 27399, 27115, 26857, 26250, 25217, 23916, 23192, 22781, 22681, 
    22890, 23328, 24176, 25289, 26513, 27164, 26925, 26176, 25684, 25220, 
    24727, 24333,
  27407, 27424, 27128, 26863, 26247, 25265, 23972, 23242, 22775, 22652, 
    22844, 23437, 24178, 25107, 26157, 27203, 26763, 26054, 25587, 25183, 
    24701, 24393,
  27193, 27214, 27113, 26863, 26293, 25254, 23979, 23194, 22804, 22657, 
    22702, 23331, 24104, 25422, 26500, 27164, 26601, 25916, 25517, 25108, 
    24714, 24219,
  26746, 26752, 27021, 26749, 26301, 25285, 24003, 23215, 22840, 22674, 
    22855, 23399, 24180, 24970, 26529, 27100, 26539, 25857, 25469, 25077, 
    24548, 24191,
  26065, 26048, 26660, 26566, 26160, 25226, 23965, 23226, 22775, 22695, 
    22964, 23432, 24153, 25114, 26343, 26794, 26589, 25974, 25579, 25164, 
    24675, 24278,
  25201, 25174, 26156, 26272, 26054, 25214, 23982, 23241, 22778, 22723, 
    22921, 23336, 24271, 25198, 26520, 26259, 26757, 26321, 25787, 25325, 
    24720, 24272,
  24281, 24262, 25583, 25924, 25906, 25248, 23948, 23209, 22813, 22683, 
    22838, 23389, 24222, 25347, 26396, 25555, 26613, 26473, 26042, 25506, 
    24892, 24359,
  23469, 23473, 25197, 25712, 25838, 25164, 23937, 23226, 22792, 22643, 
    22821, 23328, 24301, 25424, 26398, 25076, 26569, 26740, 26187, 25618, 
    24943, 24406,
  22907, 22939, 25083, 25639, 25806, 25195, 23982, 23262, 22860, 22714, 
    22904, 23391, 24104, 25237, 26816, 24967, 26819, 26782, 26284, 25704, 
    25045, 24479,
  22660, 22715, 24900, 25526, 25772, 25130, 23992, 23285, 22836, 22674, 
    22844, 23450, 24205, 25152, 26653, 24775, 26700, 26812, 26312, 25749, 
    25058, 24526,
  22701, 22752, 24789, 25426, 25660, 25125, 23951, 23288, 22839, 22717, 
    22844, 23371, 24289, 25356, 26131, 24450, 26351, 26762, 26304, 25712, 
    25064, 24426,
  22906, 22920, 24758, 25383, 25612, 25055, 23926, 23214, 22831, 22720, 
    22901, 23480, 24215, 25233, 26447, 24327, 25990, 26668, 26235, 25699, 
    25020, 24473,
  23086, 23058, 24865, 25385, 25634, 25043, 23954, 23244, 22822, 22792, 
    22875, 23417, 24239, 24998, 26459, 24335, 25890, 26631, 26249, 25754, 
    24930, 24459,
  23068, 23035, 24791, 25353, 25597, 25049, 23941, 23235, 22842, 22743, 
    22907, 23402, 24269, 25368, 26585, 24374, 25890, 26588, 26235, 25643, 
    24841, 24433,
  22791, 22787, 24626, 25243, 25531, 25046, 23930, 23229, 22804, 22766, 
    23006, 23368, 24197, 25466, 26604, 24232, 25828, 26538, 26256, 25724, 
    24975, 24359,
  22322, 22345, 24365, 25054, 25431, 24979, 23944, 23206, 22851, 22749, 
    22967, 23478, 24259, 25396, 26488, 23946, 25691, 26545, 26228, 25735, 
    25077, 24420,
  21782, 21820, 24058, 24855, 25400, 24967, 23888, 23218, 22860, 22761, 
    22938, 23422, 24210, 25161, 26450, 23673, 25635, 26545, 26318, 25681, 
    25039, 24493,
  21282, 21342, 23766, 24661, 25236, 24976, 23926, 23188, 22825, 22758, 
    23049, 23333, 24299, 25210, 26354, 23366, 25647, 26545, 26297, 25774, 
    25103, 24560,
  20901, 20996, 23650, 24640, 25194, 24917, 23902, 23242, 22898, 22784, 
    22935, 23389, 24276, 25396, 26789, 23294, 25659, 26646, 26353, 25923, 
    25199, 24574,
  20694, 20819, 23736, 24629, 25251, 24897, 23930, 23206, 22913, 22801, 
    23001, 23409, 24345, 25449, 26376, 23455, 25834, 26646, 26325, 25967, 
    25249, 24681,
  20686, 20821, 23691, 24653, 25265, 24942, 23916, 23221, 22869, 22747, 
    22899, 23432, 24215, 25254, 26498, 23483, 25834, 26632, 26326, 25874, 
    25250, 24674,
  20855, 20989, 23886, 24739, 25302, 24909, 23899, 23233, 22907, 22812, 
    22887, 23473, 24250, 25240, 26314, 23675, 25878, 26646, 26339, 26010, 
    25263, 24755,
  21145, 21276, 24190, 24939, 25365, 24889, 23854, 23251, 22840, 22792, 
    23087, 23481, 24336, 25291, 26488, 24034, 26109, 26682, 26415, 25992, 
    25314, 24789,
  21494, 21618, 24345, 24980, 25348, 24900, 23872, 23227, 22890, 22778, 
    23036, 23326, 24233, 25273, 26741, 24212, 26046, 26632, 26395, 25942, 
    25352, 24856,
  21853, 21964, 24363, 24971, 25349, 24884, 23851, 23189, 22905, 22839, 
    22967, 23364, 24144, 25278, 26307, 24125, 25816, 26545, 26340, 25935, 
    25301, 24896,
  22181, 22281, 24411, 25030, 25363, 24870, 23833, 23166, 22861, 22816, 
    23016, 23405, 24304, 25568, 26396, 24086, 25785, 26560, 26284, 25993, 
    25314, 24776,
  22461, 22541, 24523, 25139, 25343, 24853, 23827, 23151, 22805, 22828, 
    22959, 23474, 24285, 25357, 26593, 24138, 25885, 26574, 26360, 25924, 
    25276, 24876,
  22686, 22731, 24587, 25173, 25363, 24845, 23806, 23181, 22885, 22888, 
    23093, 23484, 24366, 25448, 26399, 24091, 25729, 26538, 26250, 25874, 
    25295, 24877,
  22846, 22853, 24531, 25163, 25383, 24840, 23813, 23187, 22905, 22857, 
    23094, 23451, 24216, 25634, 26581, 24054, 25698, 26539, 26271, 25812, 
    25295, 24770,
  22902, 22904, 24594, 25179, 25375, 24868, 23796, 23163, 22911, 22871, 
    23011, 23479, 24281, 25317, 26564, 24132, 25779, 26510, 26278, 25788, 
    25188, 24790,
  22814, 22847, 24579, 25204, 25395, 24784, 23768, 23202, 22853, 22777, 
    23085, 23607, 24288, 25432, 26800, 24299, 25866, 26488, 26132, 25701, 
    25137, 24750,
  22562, 22631, 24630, 25188, 25344, 24795, 23793, 23175, 22915, 22854, 
    23074, 23574, 24360, 25350, 26454, 24505, 25972, 26451, 26106, 25682, 
    25073, 24622,
  22154, 22240, 24696, 25225, 25349, 24770, 23755, 23155, 22921, 22883, 
    23008, 23500, 24360, 25609, 26846, 24675, 26172, 26337, 26029, 25570, 
    25016, 24549,
  21645, 21744, 24458, 25091, 25292, 24759, 23689, 23146, 22892, 22880, 
    23106, 23490, 24303, 25762, 26804, 24580, 26141, 26373, 26044, 25540, 
    24971, 24516,
  21157, 21304, 23979, 24808, 25206, 24672, 23727, 23129, 22933, 22910, 
    23057, 23440, 24299, 25701, 26620, 24055, 25929, 26381, 25975, 25615, 
    24927, 24456,
  20865, 21090, 23710, 24676, 25158, 24633, 23724, 23123, 22880, 22869, 
    23129, 23466, 24343, 25444, 26579, 23874, 25929, 26287, 25969, 25527, 
    24972, 24570,
  20896, 21169, 23863, 24754, 25121, 24672, 23700, 23126, 22927, 22887, 
    23066, 23565, 24247, 25491, 26506, 23926, 25910, 26388, 26051, 25640, 
    25023, 24497,
  21232, 21482, 24065, 24868, 25158, 24622, 23617, 23138, 22880, 22910, 
    23061, 23550, 24326, 25435, 26516, 24091, 25867, 26424, 26085, 25615, 
    25068, 24611,
  21723, 21910, 24388, 25027, 25213, 24614, 23648, 23159, 22925, 22899, 
    23039, 23484, 24408, 25685, 26548, 24319, 25985, 26381, 26038, 25634, 
    25113, 24571,
  22192, 22343, 24657, 25164, 25238, 24608, 23613, 23142, 22884, 22960, 
    23056, 23659, 24445, 25447, 26390, 24611, 25992, 26331, 25997, 25584, 
    25075, 24531,
  22517, 22679, 24799, 25242, 25265, 24569, 23621, 23136, 22948, 22914, 
    23113, 23652, 24408, 25593, 26907, 24789, 26129, 26324, 25990, 25616, 
    24948, 24538,
  22661, 22850, 24735, 25240, 25241, 24561, 23607, 23116, 22967, 22963, 
    23144, 23558, 24539, 25719, 26987, 24725, 26123, 26360, 26051, 25603, 
    25082, 24471,
  22666, 22863, 24660, 25186, 25193, 24550, 23607, 23172, 22952, 22958, 
    23136, 23685, 24502, 25638, 26515, 24409, 25843, 26346, 26053, 25623, 
    25107, 24512,
  22621, 22801, 24566, 25095, 25162, 24508, 23552, 23125, 22985, 22912, 
    23182, 23622, 24434, 25452, 26707, 24320, 25812, 26339, 26073, 25728, 
    25140, 24679,
  22593, 22746, 24708, 25138, 25099, 24441, 23517, 23114, 22967, 22995, 
    23097, 23661, 24527, 25659, 26754, 24467, 25993, 26325, 26067, 25691, 
    25159, 24666,
  22588, 22723, 24799, 25181, 25173, 24433, 23514, 23102, 22956, 22995, 
    23052, 23595, 24432, 25745, 26732, 24614, 26068, 26318, 26026, 25617, 
    25095, 24586,
  22585, 22721, 24840, 25273, 25145, 24396, 23521, 23087, 23029, 22981, 
    23157, 23633, 24459, 25957, 26732, 24628, 26074, 26303, 25991, 25487, 
    24981, 24513,
  22586, 22742, 24911, 25268, 25082, 24338, 23463, 23079, 22974, 22979, 
    23146, 23712, 24466, 25894, 26979, 24647, 26068, 26267, 25950, 25592, 
    24950, 24540,
  22637, 22812, 24983, 25268, 25094, 24324, 23463, 23097, 23036, 23031, 
    23186, 23636, 24614, 25954, 26973, 24722, 26193, 26310, 25950, 25580, 
    24918, 24447,
  22794, 22964, 25054, 25303, 25105, 24327, 23411, 23156, 23001, 23016, 
    23206, 23700, 24614, 25676, 26913, 24808, 26210, 26268, 25971, 25537, 
    25039, 24507,
  23077, 23216, 25170, 25354, 25017, 24238, 23387, 23101, 22957, 23034, 
    23187, 23809, 24519, 25823, 26937, 24833, 26237, 26203, 25860, 25488, 
    24880, 24307,
  23445, 23541, 25267, 25398, 25014, 24216, 23422, 23136, 22992, 23037, 
    23241, 23685, 24704, 25816, 26932, 24928, 26256, 26160, 25813, 25388, 
    24798, 24347,
  23822, 23872, 25396, 25409, 24997, 24176, 23356, 23086, 23028, 23049, 
    23284, 23711, 24652, 26060, 27114, 24902, 26181, 26124, 25765, 25382, 
    24741, 24247,
  24152, 24149, 25401, 25403, 24981, 24143, 23370, 23096, 23046, 23064, 
    23242, 23779, 24615, 26034, 27029, 24642, 25864, 26067, 25751, 25314, 
    24792, 24381,
  24400, 24338, 25376, 25390, 24858, 24071, 23339, 23084, 23060, 23055, 
    23179, 23843, 24771, 25809, 26832, 24237, 25690, 26117, 25793, 25396, 
    24901, 24502,
  24497, 24388, 25288, 25322, 24866, 24031, 23297, 23102, 23055, 23084, 
    23276, 23816, 24690, 26010, 27382, 23933, 25634, 26088, 25751, 25396, 
    24831, 24482,
  24379, 24250, 25260, 25245, 24758, 23970, 23309, 23114, 23055, 23084, 
    23405, 23890, 24825, 26137, 27168, 23656, 25429, 25966, 25622, 25197, 
    24787, 24322,
  24136, 24005, 25260, 25191, 24721, 23886, 23267, 23087, 23070, 23125, 
    23356, 23880, 24821, 26023, 27243, 23731, 25447, 25829, 25505, 25117, 
    24628, 24242,
  24009, 23880, 25260, 25170, 24655, 23822, 23243, 23117, 23050, 23085, 
    23303, 23959, 24853, 26290, 27204, 24001, 25703, 25685, 25402, 24999, 
    24482, 24008 ;
}
