netcdf icec_mirs_snpp_1 {
dimensions:
	Scanline = 12 ;
	Field_of_view = 96 ;
	Channel = 22 ;
	Qc_dim = 4 ;
variables:
	short Atm_type(Scanline, Field_of_view) ;
		Atm_type:description = "type of atmosphere:currently missing" ;
		Atm_type:coordinates = "Longitude Latitude" ;
	short BT(Scanline, Field_of_view, Channel) ;
		BT:long_name = "Channel Temperature (K)" ;
		BT:units = "Kelvin" ;
		BT:coordinates = "Longitude Latitude Freq" ;
		BT:scale_factor = 0.01 ;
		BT:_FillValue = -999s ;
		BT:valid_range = 0, 50000 ;
	short CLW(Scanline, Field_of_view) ;
		CLW:long_name = "Cloud liquid Water (mm)" ;
		CLW:units = "mm" ;
		CLW:coordinates = "Longitude Latitude" ;
		CLW:scale_factor = 0.01 ;
		CLW:_FillValue = -999s ;
		CLW:valid_range = 0, 10000 ;
	short ChanSel(Scanline, Field_of_view, Channel) ;
		ChanSel:long_name = "Channels Selection Used in Retrieval" ;
		ChanSel:units = "1" ;
		ChanSel:coordinates = "Longitude Latitude Freq" ;
		ChanSel:_FillValue = -999s ;
		ChanSel:valid_range = 0, 1 ;
	float ChiSqr(Scanline, Field_of_view) ;
		ChiSqr:description = "Convergence rate: <3-good,>10-bad" ;
		ChiSqr:units = "1" ;
		ChiSqr:coordinates = "Longitude Latitude" ;
		ChiSqr:_FillValue = -999.f ;
		ChiSqr:valid_range = 0.f, 1000.f ;
	short CldBase(Scanline, Field_of_view) ;
		CldBase:long_name = "Cloud Base Pressure" ;
		CldBase:scale_factor = 0.1 ;
		CldBase:coordinates = "Longitude Latitude" ;
	short CldThick(Scanline, Field_of_view) ;
		CldThick:long_name = "Cloud Thickness" ;
		CldThick:scale_factor = 0.1 ;
		CldThick:coordinates = "Longitude Latitude" ;
	short CldTop(Scanline, Field_of_view) ;
		CldTop:long_name = "Cloud Top Pressure" ;
		CldTop:scale_factor = 0.1 ;
		CldTop:coordinates = "Longitude Latitude" ;
	short Emis(Scanline, Field_of_view, Channel) ;
		Emis:long_name = "Channel Emissivity" ;
		Emis:units = "1" ;
		Emis:coordinates = "Longitude Latitude Freq" ;
		Emis:scale_factor = 0.0001 ;
		Emis:_FillValue = -999s ;
		Emis:valid_range = 0, 10000 ;
	float Freq(Channel) ;
		Freq:description = "Central Frequencies (GHz)" ;
	short GWP(Scanline, Field_of_view) ;
		GWP:long_name = "Graupel Water Path (mm)" ;
		GWP:units = "mm" ;
		GWP:coordinates = "Longitude Latitude" ;
		GWP:scale_factor = 0.01 ;
		GWP:_FillValue = -999s ;
		GWP:valid_range = 0, 10000 ;
	short IWP(Scanline, Field_of_view) ;
		IWP:long_name = "Ice Water Path (mm)" ;
		IWP:units = "mm" ;
		IWP:coordinates = "Longitude Latitude" ;
		IWP:scale_factor = 0.01 ;
		IWP:_FillValue = -999s ;
		IWP:valid_range = 0, 10000 ;
	short LWP(Scanline, Field_of_view) ;
		LWP:long_name = "Liquid Water Path (mm)" ;
		LWP:units = "mm" ;
		LWP:coordinates = "Longitude Latitude" ;
		LWP:scale_factor = 0.01 ;
		LWP:_FillValue = -999s ;
		LWP:valid_range = 0, 10000 ;
	float LZ_angle(Scanline, Field_of_view) ;
		LZ_angle:long_name = "Local Zenith Angle degree" ;
		LZ_angle:units = "degrees" ;
		LZ_angle:coordinates = "Longitude Latitude" ;
		LZ_angle:_FillValue = -999.f ;
		LZ_angle:valid_range = -70.f, 70.f ;
	float Latitude(Scanline, Field_of_view) ;
		Latitude:long_name = "Latitude of the view (-90,90)" ;
		Latitude:units = "degrees" ;
		Latitude:_FillValue = -999.f ;
		Latitude:valid_range = -90.f, 90.f ;
	float Longitude(Scanline, Field_of_view) ;
		Longitude:long_name = "Longitude of the view (-180,180)" ;
		Longitude:units = "degrees" ;
		Longitude:_FillValue = -999.f ;
		Longitude:valid_range = -180.f, 180.f ;
	short Orb_mode(Scanline) ;
		Orb_mode:description = "0-ascending,1-descending" ;
		Orb_mode:units = "1" ;
		Orb_mode:_FillValue = -999s ;
		Orb_mode:valid_range = 0, 1 ;
	short Polo(Channel) ;
		Polo:description = "Polarizations" ;
	short PrecipType(Scanline, Field_of_view) ;
		PrecipType:long_name = "Precipitation Type (Frozen/Liquid)" ;
		PrecipType:coordinates = "Longitude Latitude" ;
	short Prob_SF(Scanline, Field_of_view) ;
		Prob_SF:long_name = "Probability of falling snow (%)" ;
		Prob_SF:units = "percent" ;
		Prob_SF:coordinates = "Longitude Latitude" ;
		Prob_SF:_FillValue = -999s ;
		Prob_SF:valid_range = 0, 100 ;
	short Qc(Scanline, Field_of_view, Qc_dim) ;
		Qc:description = "Qc: 0-good, 1-usable with problem, 2-bad" ;
	float RAzi_angle(Scanline, Field_of_view) ;
		RAzi_angle:long_name = "Relative Azimuth Angle 0-360 degree" ;
		RAzi_angle:coordinates = "Longitude Latitude" ;
	short RFlag(Scanline, Field_of_view) ;
		RFlag:long_name = "Rain Flag" ;
		RFlag:coordinates = "Longitude Latitude" ;
	short RR(Scanline, Field_of_view) ;
		RR:long_name = "Rain Rate (mm/hr)" ;
		RR:units = "mm/hr" ;
		RR:coordinates = "Longitude Latitude" ;
		RR:scale_factor = 0.1 ;
		RR:_FillValue = -999s ;
		RR:valid_range = 0, 1000 ;
	short RWP(Scanline, Field_of_view) ;
		RWP:long_name = "Rain Water Path (mm)" ;
		RWP:units = "mm" ;
		RWP:coordinates = "Longitude Latitude" ;
		RWP:scale_factor = 0.01 ;
		RWP:_FillValue = -999s ;
		RWP:valid_range = 0, 10000 ;
	short SFR(Scanline, Field_of_view) ;
		SFR:long_name = "Snow Fall Rate in mm/hr" ;
		SFR:units = "mm/hr" ;
		SFR:coordinates = "Longitude Latitude" ;
		SFR:scale_factor = 0.01 ;
		SFR:_FillValue = -999s ;
		SFR:valid_range = 0, 10000 ;
	short SIce(Scanline, Field_of_view) ;
		SIce:long_name = "Sea Ice Concentration (%)" ;
		SIce:units = "percent" ;
		SIce:coordinates = "Longitude Latitude" ;
		SIce:_FillValue = -999s ;
		SIce:valid_range = 0, 100 ;
	short SIce_FY(Scanline, Field_of_view) ;
		SIce_FY:long_name = "First-Year Sea Ice Concentration (%)" ;
		SIce_FY:units = "percent" ;
		SIce_FY:coordinates = "Longitude Latitude" ;
		SIce_FY:_FillValue = -999s ;
		SIce_FY:valid_range = 0, 100 ;
	short SIce_MY(Scanline, Field_of_view) ;
		SIce_MY:long_name = "Multi-Year Sea Ice Concentration (%)" ;
		SIce_MY:units = "percent" ;
		SIce_MY:coordinates = "Longitude Latitude" ;
		SIce_MY:_FillValue = -999s ;
		SIce_MY:valid_range = 0, 100 ;
	short SWE(Scanline, Field_of_view) ;
		SWE:long_name = "Snow Water Equivalent (cm)" ;
		SWE:units = "cm" ;
		SWE:coordinates = "Longitude Latitude" ;
		SWE:scale_factor = 0.01 ;
		SWE:_FillValue = -999s ;
		SWE:valid_range = 0, 10000 ;
	short SWP(Scanline, Field_of_view) ;
		SWP:long_name = "Snow Water Path" ;
		SWP:units = "mm" ;
		SWP:coordinates = "Longitude Latitude" ;
		SWP:scale_factor = 0.01 ;
		SWP:_FillValue = -999s ;
		SWP:valid_range = 0, 10000 ;
	float SZ_angle(Scanline, Field_of_view) ;
		SZ_angle:long_name = "Solar Zenith Angle (-90,90) degree" ;
		SZ_angle:coordinates = "Longitude Latitude" ;
	double ScanTime_UTC(Scanline) ;
		ScanTime_UTC:long_name = "Number of seconds since 00:00:00 UTC" ;
		ScanTime_UTC:units = "seconds" ;
		ScanTime_UTC:_FillValue = -999. ;
		ScanTime_UTC:valid_range = 0., 86400. ;
	short ScanTime_dom(Scanline) ;
		ScanTime_dom:long_name = "Calendar day of the month 1-31" ;
		ScanTime_dom:units = "days" ;
		ScanTime_dom:_FillValue = -999s ;
		ScanTime_dom:valid_range = 1, 31 ;
	short ScanTime_doy(Scanline) ;
		ScanTime_doy:long_name = "julian day 1-366" ;
		ScanTime_doy:units = "days" ;
		ScanTime_doy:_FillValue = -999s ;
		ScanTime_doy:valid_range = 1, 366 ;
	short ScanTime_hour(Scanline) ;
		ScanTime_hour:long_name = "hour of the day 0-23" ;
		ScanTime_hour:units = "hours" ;
		ScanTime_hour:_FillValue = -999s ;
		ScanTime_hour:valid_range = 0, 23 ;
	short ScanTime_minute(Scanline) ;
		ScanTime_minute:long_name = "minute of the hour 0-59" ;
		ScanTime_minute:units = "minutes" ;
		ScanTime_minute:_FillValue = -999s ;
		ScanTime_minute:valid_range = 0, 59 ;
	short ScanTime_month(Scanline) ;
		ScanTime_month:long_name = "Calendar month 1-12" ;
		ScanTime_month:units = "months" ;
		ScanTime_month:_FillValue = -999s ;
		ScanTime_month:valid_range = 1, 12 ;
	short ScanTime_second(Scanline) ;
		ScanTime_second:long_name = "second of the minute 0-59" ;
		ScanTime_second:units = "seconds" ;
		ScanTime_second:_FillValue = -999s ;
		ScanTime_second:valid_range = 0, 59 ;
	short ScanTime_year(Scanline) ;
		ScanTime_year:long_name = "Calendar Year 20XX" ;
		ScanTime_year:units = "years" ;
		ScanTime_year:_FillValue = -999s ;
		ScanTime_year:valid_range = 2011, 2050 ;
	short Sfc_type(Scanline, Field_of_view) ;
		Sfc_type:description = "type of surface:0-ocean,1-sea ice,2-land,3-snow" ;
		Sfc_type:units = "1" ;
		Sfc_type:coordinates = "Longitude Latitude" ;
		Sfc_type:_FillValue = -999s ;
		Sfc_type:valid_range = 0, 3 ;
	short Snow(Scanline, Field_of_view) ;
		Snow:long_name = "Snow Cover" ;
		Snow:units = "1" ;
		Snow:coordinates = "Longitude Latitude" ;
		Snow:_FillValue = -999s ;
		Snow:valid_range = 0, 1 ;
	short SnowGS(Scanline, Field_of_view) ;
		SnowGS:long_name = "Snow Grain Size (mm)" ;
		SnowGS:units = "mm" ;
		SnowGS:coordinates = "Longitude Latitude" ;
		SnowGS:scale_factor = 0.01 ;
		SnowGS:_FillValue = -999s ;
		SnowGS:valid_range = 0, 2000 ;
	short SurfM(Scanline, Field_of_view) ;
		SurfM:long_name = "Surface Moisture" ;
		SurfM:scale_factor = 0.1 ;
		SurfM:coordinates = "Longitude Latitude" ;
	short SurfP(Scanline, Field_of_view) ;
		SurfP:long_name = "Surface Pressure (mb)" ;
		SurfP:units = "millibars" ;
		SurfP:coordinates = "Longitude Latitude" ;
		SurfP:scale_factor = 0.1 ;
		SurfP:_FillValue = -999s ;
		SurfP:valid_range = 0, 12000 ;
	short TPW(Scanline, Field_of_view) ;
		TPW:long_name = "Total Precipitable Water (mm)" ;
		TPW:units = "mm" ;
		TPW:coordinates = "Longitude Latitude" ;
		TPW:scale_factor = 0.1 ;
		TPW:_FillValue = -999s ;
		TPW:valid_range = 0, 2000 ;
	short TSkin(Scanline, Field_of_view) ;
		TSkin:long_name = "Skin Temperature (K)" ;
		TSkin:units = "Kelvin" ;
		TSkin:coordinates = "Longitude Latitude" ;
		TSkin:scale_factor = 0.01 ;
		TSkin:_FillValue = -999s ;
		TSkin:valid_range = 0, 40000 ;
	short WindDir(Scanline, Field_of_view) ;
		WindDir:long_name = "Wind Direction" ;
		WindDir:scale_factor = 0.01 ;
		WindDir:coordinates = "Longitude Latitude" ;
	short WindSp(Scanline, Field_of_view) ;
		WindSp:long_name = "Wind Speed (m/s)" ;
		WindSp:scale_factor = 0.01 ;
		WindSp:coordinates = "Longitude Latitude" ;
	short WindU(Scanline, Field_of_view) ;
		WindU:long_name = "U-direction Wind Speed (m/s)" ;
		WindU:scale_factor = 0.01 ;
		WindU:coordinates = "Longitude Latitude" ;
	short WindV(Scanline, Field_of_view) ;
		WindV:long_name = "V-direction Wind Speed (m/s)" ;
		WindV:scale_factor = 0.01 ;
		WindV:coordinates = "Longitude Latitude" ;
	short YM(Scanline, Field_of_view, Channel) ;
		YM:long_name = "Un-Corrected Channel Temperature (K)" ;
		YM:units = "Kelvin" ;
		YM:coordinates = "Longitude Latitude Freq" ;
		YM:scale_factor = 0.01 ;
		YM:_FillValue = -999s ;
		YM:valid_range = 0, 50000 ;

// global attributes:
		:missing_value = -999 ;
		:notretrievedproduct_value = -888 ;
		:noretrieval_value = -99 ;
		:cdf_version = 4. ;
		:alg_version = 4201 ;
		:dap_version = "v11r4" ;
		:Conventions = "CF-1.5" ;
		:Metadata_Conventions = "CF-1.5, Unidata Dataset Discovery v1.0" ;
		:standard_name_vocabulary = "CF Standard Name Table (version 17, 24 March 2011)" ;
		:project = "Microwave Integrated Retrieval System" ;
		:title = "MIRS IMG" ;
		:summary = "MIRS imaging products including surface emissivity, TPW, CLW, RWP, IWP, LST." ;
		:date_created = "2021-06-30T02:01:08Z" ;
		:institution = "DOC/NOAA/NESDIS/NDE > NPOESS Data Exploitation, NESDIS, NOAA, U.S. Department of Commerce" ;
		:naming_authority = "gov.noaa.nesdis.nde" ;
		:production_site = "NSOF" ;
		:production_environment = "OE" ;
		:satellite_name = "NPP" ;
		:instrument_name = "ATMS" ;
		:creator_name = "DOC/NOAA/NESDIS/STAR > MIRS TEAM, Center for Satellite Applications and Research, NESDIS, NOAA, U.S. Department of Commerce" ;
		:creator_email = "Christopher.Grassotti@noaa.gov, Quanhua.Liu@noaa.gov, Shu-yan.Liu@noaa.gov, ryan.honeyager@noaa.gov, Yong-Keun.Lee@noaa.gov " ;
		:creator_url = "http://www.star.nesdis.noaa.gov/mirs" ;
		:publisher_name = "DOC/NOAA/NESDIS/NDE > NPOESS Data Exploitation, NESDIS, NOAA, U.S. Department of Commerce" ;
		:publisher_email = "NDE_POC@noaa.gov" ;
		:publisher_url = "http://projects.osd.noaa.gov/NDE" ;
		:Metadata_Link = "NDE product-specific output file name" ;
		:references = "http://www.star.nesdis.noaa.gov/mirs/documentation.php" ;
		:history = "Mon Jul 29 20:07:53 2024: ncks NPR-MIRS-IMG_v11r4_npp_s202106300127066_e202106300127383_c202106300201000.nc icec_mirs_snpp_1.nc\nCreated by MIRS Version 11.4" ;
		:processing_level = "NOAA Level 2 data" ;
		:source = "SATMS_npp_d20210630_t0127066_e0127383_b50120_c20210630015713485030_oebc_ops.h5" ;
		:time_coverage_start = "2021-06-30T01:27:06Z" ;
		:time_coverage_end = "2021-06-30T01:27:38Z" ;
		:cdm_data_type = "Swath" ;
		:geospatial_lat_units = "degrees_north" ;
		:geospatial_lon_units = "degrees_east" ;
		:geospatial_lat_resolution = "100" ;
		:geospatial_lon_resolution = "100" ;
		:geospatial_first_scanline_first_fov_lat = 61.18f ;
		:geospatial_first_scanline_first_fov_lon = 135.75f ;
		:geospatial_first_scanline_last_fov_lat = 69.42f ;
		:geospatial_first_scanline_last_fov_lon = -171.14f ;
		:geospatial_last_scanline_first_fov_lat = 62.38f ;
		:geospatial_last_scanline_first_fov_lon = 133.09f ;
		:geospatial_last_scanline_last_fov_lat = 71.1f ;
		:geospatial_last_scanline_last_fov_lon = -170.7f ;
		:total_number_retrievals = 1152 ;
		:percentage_optimal_retrievals = 0.3125f ;
		:percentage_suboptimal_retrievals = 0.6875f ;
		:percentage_bad_retrievals = 0.f ;
		:start_orbit_number = 50120 ;
		:end_orbit_number = 50120 ;
		:id = "ndepgsl-op-13_2021-06-30T02:01:08Z_0000001764860342_SATMS_npp_d20210630_t0127066_e0127383_b50120_c20210630015713485030_oebc_ops.h5" ;
		:NCO = "netCDF Operators version 5.0.6 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco)" ;
data:

 Atm_type =
  -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999,
  -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999,
  -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999,
  -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999,
  -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999,
  -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999,
  -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999,
  -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999,
  -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999,
  -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999,
  -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999,
  -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, 
    -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999, -999 ;

 BT =
  28033, 28007, 27902, 27183, 25827, 24165, 22717, 22271, 22167, 22482, 
    22861, 23661, 24690, 25965, 26442, 28537, 28843, 28000, 27396, 26801, 
    26001, 25170,
  28028, 28003, 27960, 27247, 25997, 24305, 22803, 22294, 22167, 22530, 
    22834, 23621, 24794, 25776, 26497, 28554, 28913, 27954, 27369, 26851, 
    25989, 25016,
  28005, 28003, 27832, 27312, 26097, 24389, 22935, 22362, 22200, 22486, 
    22914, 23612, 24536, 25778, 26890, 28420, 28719, 27964, 27309, 26807, 
    26016, 25017,
  27927, 27971, 27810, 27310, 26166, 24501, 22948, 22366, 22168, 22519, 
    22904, 23552, 24540, 25775, 26588, 28251, 28670, 27847, 27249, 26689, 
    25996, 24996,
  27886, 27966, 27741, 27339, 26255, 24612, 23047, 22352, 22206, 22547, 
    22929, 23512, 24465, 25796, 26509, 28179, 28601, 27816, 27153, 26552, 
    25806, 24922,
  27875, 27983, 27735, 27337, 26341, 24704, 23095, 22472, 22247, 22501, 
    22862, 23540, 24592, 25667, 26685, 28139, 28562, 27767, 27148, 26478, 
    25660, 24774,
  27914, 28025, 27763, 27424, 26437, 24843, 23165, 22472, 22214, 22479, 
    22875, 23503, 24474, 25573, 26453, 28338, 28706, 27879, 27119, 26478, 
    25616, 24681,
  27999, 28103, 27949, 27547, 26589, 24887, 23226, 22520, 22237, 22488, 
    22865, 23523, 24483, 25700, 26359, 28432, 28916, 27921, 27186, 26422, 
    25552, 24687,
  28085, 28185, 27986, 27628, 26649, 25000, 23312, 22569, 22229, 22448, 
    22868, 23462, 24481, 25601, 26503, 28499, 28916, 27859, 27121, 26478, 
    25495, 24540,
  28109, 28220, 28018, 27657, 26697, 25050, 23387, 22610, 22268, 22456, 
    22871, 23490, 24488, 25569, 26556, 28474, 28835, 27856, 27028, 26323, 
    25291, 24293,
  28066, 28191, 27925, 27633, 26687, 25093, 23434, 22651, 22269, 22430, 
    22804, 23489, 24420, 25510, 26447, 28422, 28849, 27675, 26896, 26091, 
    25042, 24190,
  27999, 28134, 27778, 27516, 26632, 25087, 23465, 22673, 22272, 22438, 
    22992, 23424, 24419, 25495, 26492, 28245, 28522, 27506, 26756, 25859, 
    24984, 24057,
  27917, 28058, 27676, 27487, 26687, 25207, 23522, 22723, 22298, 22486, 
    22910, 23421, 24364, 25376, 26660, 28048, 28340, 27500, 26656, 25837, 
    24790, 24022,
  27819, 27949, 27704, 27480, 26726, 25241, 23554, 22733, 22341, 22534, 
    22890, 23469, 24610, 25616, 26153, 28077, 28511, 27582, 26769, 25928, 
    24884, 24066,
  27697, 27829, 27628, 27444, 26725, 25301, 23650, 22762, 22305, 22436, 
    22954, 23407, 24364, 25601, 26500, 28044, 28497, 27631, 26835, 26038, 
    24938, 24082,
  27588, 27732, 27501, 27369, 26704, 25330, 23635, 22802, 22361, 22482, 
    22822, 23402, 24351, 25440, 26674, 27849, 28384, 27679, 26924, 26028, 
    25096, 24260,
  27520, 27682, 27394, 27223, 26708, 25314, 23687, 22845, 22386, 22507, 
    22857, 23469, 24273, 25515, 26622, 27687, 28309, 27574, 26744, 25896, 
    24953, 24239,
  27510, 27675, 27323, 27263, 26728, 25390, 23729, 22836, 22368, 22471, 
    22851, 23483, 24207, 25534, 26444, 27673, 28321, 27384, 26537, 25704, 
    24914, 24150,
  27535, 27700, 27436, 27335, 26772, 25432, 23791, 22876, 22382, 22470, 
    22806, 23353, 24419, 25250, 26328, 27793, 28323, 27254, 26426, 25684, 
    24887, 24256,
  27579, 27744, 27484, 27354, 26802, 25470, 23805, 22926, 22440, 22434, 
    22874, 23358, 24245, 25499, 26535, 27841, 28141, 27002, 26191, 25509, 
    24900, 24316,
  27619, 27803, 27556, 27376, 26830, 25507, 23830, 22919, 22410, 22499, 
    22767, 23344, 24411, 25507, 26656, 27853, 28118, 26951, 26200, 25436, 
    24746, 24115,
  27663, 27861, 27532, 27382, 26829, 25537, 23850, 22951, 22473, 22495, 
    22825, 23382, 24336, 25389, 26625, 27943, 28176, 26943, 26124, 25411, 
    24810, 24128,
  27707, 27892, 27481, 27307, 26806, 25541, 23895, 23018, 22437, 22429, 
    22807, 23365, 24218, 25378, 26414, 27888, 28049, 26872, 26147, 25479, 
    24778, 24134,
  27701, 27845, 27399, 27299, 26763, 25528, 23904, 23010, 22481, 22415, 
    22853, 23393, 24381, 25475, 26712, 27770, 27821, 26810, 26210, 25559, 
    24860, 24260,
  27571, 27647, 27434, 27273, 26725, 25543, 23946, 23001, 22507, 22479, 
    22756, 23262, 24239, 25391, 26512, 27838, 27820, 26771, 26153, 25539, 
    24826, 24237,
  27291, 27292, 27382, 27212, 26753, 25557, 23948, 23049, 22498, 22426, 
    22765, 23299, 24172, 25184, 26399, 27826, 27829, 26688, 26050, 25512, 
    24856, 24115,
  26933, 26878, 27053, 27074, 26671, 25522, 23976, 23044, 22518, 22455, 
    22865, 23366, 24210, 25531, 26264, 27528, 27701, 26696, 26026, 25454, 
    24751, 24194,
  26643, 26568, 26722, 26853, 26592, 25478, 23982, 23073, 22506, 22463, 
    22659, 23271, 24257, 25387, 26044, 27185, 27663, 26630, 26037, 25496, 
    24790, 24212,
  26547, 26466, 26504, 26710, 26544, 25506, 23994, 23086, 22514, 22503, 
    22783, 23321, 24170, 25320, 26293, 27030, 27472, 26566, 26020, 25482, 
    24763, 24099,
  26669, 26584, 26704, 26851, 26572, 25571, 24010, 23071, 22581, 22514, 
    22786, 23299, 24009, 25538, 26348, 27140, 27513, 26549, 25975, 25443, 
    24724, 24112,
  26914, 26844, 26991, 27017, 26657, 25569, 24039, 23136, 22577, 22526, 
    22864, 23354, 24276, 25259, 26387, 27409, 27673, 26609, 25959, 25454, 
    24737, 24141,
  27150, 27138, 27085, 27103, 26714, 25587, 24029, 23149, 22557, 22506, 
    22791, 23318, 24161, 25229, 26595, 27585, 27729, 26563, 25916, 25311, 
    24744, 24181,
  27297, 27355, 27128, 27119, 26698, 25609, 24055, 23125, 22605, 22517, 
    22793, 23388, 24287, 25417, 26410, 27585, 27798, 26488, 25901, 25310, 
    24763, 24134,
  27363, 27444, 27269, 27198, 26741, 25629, 24097, 23139, 22628, 22561, 
    22775, 23359, 24132, 25375, 26435, 27621, 27681, 26487, 25913, 25361, 
    24686, 24121,
  27380, 27446, 27356, 27193, 26720, 25603, 24058, 23142, 22608, 22580, 
    22829, 23404, 24213, 25392, 26363, 27737, 27570, 26484, 25907, 25294, 
    24660, 24161,
  27362, 27421, 27373, 27188, 26762, 25574, 24065, 23174, 22601, 22527, 
    22856, 23378, 24161, 25331, 26366, 27685, 27534, 26490, 25844, 25344, 
    24691, 24066,
  27310, 27398, 27288, 27102, 26691, 25592, 24092, 23177, 22623, 22495, 
    22737, 23239, 24249, 25457, 26719, 27567, 27445, 26467, 25810, 25343, 
    24717, 24270,
  27234, 27350, 27135, 27011, 26575, 25578, 24095, 23183, 22664, 22504, 
    22779, 23208, 24181, 25367, 26154, 27388, 27213, 26387, 25824, 25392, 
    24755, 24183,
  27144, 27275, 26913, 26838, 26500, 25510, 24104, 23219, 22682, 22554, 
    22852, 23395, 24193, 25313, 26128, 27108, 26878, 26115, 25686, 25224, 
    24653, 24171,
  27049, 27178, 26771, 26690, 26384, 25473, 24088, 23194, 22675, 22547, 
    22818, 23413, 24203, 25360, 26444, 26857, 26404, 25944, 25534, 25199, 
    24615, 24085,
  26947, 27067, 26652, 26632, 26278, 25443, 24108, 23218, 22685, 22558, 
    22800, 23295, 24244, 25411, 26450, 26738, 26241, 25993, 25643, 25310, 
    24679, 24212,
  26838, 26937, 26576, 26507, 26250, 25390, 24031, 23204, 22651, 22621, 
    22824, 23310, 24110, 25363, 26579, 26661, 26456, 26166, 25801, 25310, 
    24719, 24128,
  26738, 26809, 26526, 26504, 26207, 25379, 24054, 23223, 22655, 22610, 
    22873, 23397, 24157, 25289, 26453, 26525, 26446, 26140, 25773, 25375, 
    24726, 24203,
  26681, 26722, 26469, 26463, 26209, 25379, 24070, 23215, 22647, 22590, 
    22792, 23317, 24312, 25526, 26725, 26488, 26304, 26174, 25776, 25287, 
    24701, 24276,
  26686, 26718, 26553, 26569, 26262, 25437, 24073, 23253, 22682, 22536, 
    22926, 23292, 24305, 25349, 26371, 26532, 26518, 26274, 25822, 25331, 
    24763, 24176,
  26755, 26795, 26693, 26636, 26304, 25404, 24132, 23231, 22744, 22582, 
    22834, 23311, 24229, 25355, 26708, 26618, 26662, 26317, 25916, 25369, 
    24745, 24203,
  26832, 26887, 26751, 26709, 26367, 25437, 24151, 23274, 22707, 22570, 
    22912, 23332, 24199, 25314, 26515, 26708, 26824, 26401, 25990, 25415, 
    24866, 24261,
  26874, 26938, 26731, 26759, 26373, 25509, 24156, 23220, 22716, 22625, 
    22870, 23385, 24376, 25389, 26165, 26823, 26969, 26432, 25985, 25447, 
    24864, 24365,
  26864, 26950, 26737, 26716, 26361, 25467, 24104, 23272, 22739, 22701, 
    22884, 23438, 24206, 25549, 26385, 26787, 26860, 26365, 25899, 25474, 
    24844, 24278,
  26844, 26958, 26685, 26681, 26330, 25376, 24093, 23317, 22707, 22627, 
    22801, 23319, 24251, 25418, 26598, 26610, 26591, 26247, 25821, 25348, 
    24851, 24264,
  26840, 26971, 26623, 26575, 26287, 25464, 24110, 23236, 22739, 22584, 
    22876, 23408, 24232, 25511, 26573, 26557, 26747, 26335, 25887, 25400, 
    24749, 24244,
  26862, 26976, 26707, 26661, 26351, 25467, 24116, 23269, 22753, 22707, 
    22889, 23334, 24169, 25404, 26372, 26616, 26721, 26388, 25871, 25366, 
    24716, 24090,
  26856, 26941, 26820, 26760, 26374, 25464, 24055, 23234, 22690, 22620, 
    22896, 23446, 24245, 25385, 26629, 26768, 26816, 26340, 25880, 25374, 
    24666, 24278,
  26748, 26806, 26835, 26812, 26400, 25444, 24102, 23279, 22724, 22666, 
    22880, 23382, 24287, 25314, 26215, 26888, 26737, 26356, 25869, 25295, 
    24724, 24097,
  26498, 26553, 26756, 26726, 26350, 25431, 24065, 23265, 22757, 22650, 
    22871, 23308, 24164, 25328, 26488, 26816, 26544, 26169, 25752, 25302, 
    24774, 24138,
  26146, 26225, 26489, 26523, 26289, 25401, 24130, 23283, 22751, 22694, 
    22983, 23362, 24259, 25380, 26246, 26550, 26071, 25768, 25631, 25159, 
    24647, 24125,
  25830, 25944, 26169, 26410, 26282, 25420, 24069, 23260, 22785, 22710, 
    22867, 23352, 24286, 25450, 26799, 26278, 25878, 25681, 25512, 25135, 
    24641, 24212,
  25723, 25842, 26212, 26356, 26219, 25396, 24083, 23242, 22812, 22647, 
    22825, 23390, 24276, 25315, 25942, 26244, 26415, 25966, 25588, 25160, 
    24622, 24119,
  25908, 26019, 26338, 26496, 26302, 25356, 24057, 23264, 22792, 22670, 
    22973, 23460, 24335, 25432, 26634, 26496, 26762, 26202, 25692, 25247, 
    24661, 24072,
  26317, 26439, 26763, 26772, 26437, 25440, 24038, 23258, 22779, 22671, 
    22841, 23401, 24106, 25354, 26354, 27037, 27309, 26445, 25828, 25342, 
    24733, 24153,
  26800, 26967, 27174, 27019, 26512, 25482, 24073, 23235, 22806, 22723, 
    23001, 23389, 24290, 25362, 26629, 27453, 27611, 26507, 25853, 25285, 
    24684, 24107,
  27187, 27417, 27259, 27066, 26556, 25452, 24053, 23280, 22762, 22725, 
    22979, 23340, 24229, 25478, 26259, 27628, 27708, 26621, 25938, 25293, 
    24685, 24034,
  27401, 27665, 27255, 27046, 26532, 25378, 24012, 23207, 22756, 22691, 
    22834, 23278, 24267, 25271, 26732, 27586, 27646, 26684, 25974, 25331, 
    24667, 24126,
  27474, 27710, 27187, 27021, 26543, 25424, 24036, 23234, 22791, 22742, 
    22903, 23311, 24326, 25327, 26547, 27523, 27733, 26732, 26049, 25343, 
    24668, 23993,
  27461, 27649, 27197, 26976, 26471, 25383, 24009, 23244, 22797, 22692, 
    22894, 23443, 24354, 25380, 26320, 27513, 27646, 26790, 26071, 25387, 
    24751, 24221,
  27404, 27562, 27177, 27013, 26484, 25407, 23950, 23237, 22795, 22751, 
    22985, 23434, 24213, 25410, 26625, 27476, 27582, 26781, 26094, 25418, 
    24643, 24201,
  27326, 27495, 27104, 26966, 26512, 25375, 23987, 23203, 22768, 22712, 
    22964, 23377, 24152, 25365, 26644, 27421, 27575, 26774, 26056, 25336, 
    24765, 24201,
  27236, 27451, 27024, 26926, 26405, 25323, 23946, 23199, 22758, 22776, 
    22965, 23533, 24415, 25411, 26554, 27329, 27612, 26813, 26104, 25387, 
    24689, 24144,
  27168, 27421, 26872, 26866, 26404, 25275, 23904, 23155, 22800, 22699, 
    22973, 23376, 24163, 25512, 26800, 27205, 27540, 26807, 26145, 25404, 
    24741, 24105,
  27158, 27396, 26818, 26788, 26270, 25250, 23847, 23154, 22779, 22740, 
    22962, 23497, 24266, 25521, 26645, 27096, 27401, 26797, 26197, 25412, 
    24717, 24166,
  27159, 27337, 26779, 26759, 26255, 25156, 23849, 23190, 22768, 22770, 
    22933, 23426, 24387, 25440, 26826, 27068, 27387, 26765, 26066, 25366, 
    24676, 24040,
  27002, 27102, 26775, 26673, 26203, 25175, 23881, 23157, 22772, 22804, 
    22963, 23423, 24449, 25494, 26805, 27068, 27192, 26510, 25972, 25276, 
    24561, 24132,
  26408, 26454, 26832, 26743, 26220, 25113, 23823, 23140, 22800, 22833, 
    22989, 23508, 24323, 25558, 26795, 27082, 27376, 26754, 26233, 25557, 
    24850, 24234,
  25203, 25231, 26655, 26619, 26175, 25113, 23823, 23171, 22798, 22832, 
    23065, 23445, 24300, 25653, 26409, 27035, 27548, 26967, 26335, 25623, 
    24845, 24161,
  23541, 23619, 25654, 26015, 25956, 25029, 23726, 23126, 22790, 22778, 
    23011, 23506, 24260, 25434, 26705, 26246, 27434, 26935, 26342, 25694, 
    24898, 24209,
  22007, 22186, 23805, 24968, 25517, 24907, 23725, 23137, 22862, 22787, 
    23012, 23426, 24405, 25593, 26787, 24051, 26258, 26833, 26411, 25806, 
    25012, 24359,
  21297, 21594, 22657, 24326, 25271, 24827, 23711, 23147, 22793, 22814, 
    23063, 23531, 24464, 25741, 26400, 22306, 25146, 26687, 26411, 25872, 
    25186, 24437,
  21792, 22110, 23348, 24717, 25373, 24835, 23709, 23083, 22809, 22836, 
    23124, 23587, 24365, 25694, 26819, 22955, 25377, 26763, 26457, 25973, 
    25219, 24553,
  23203, 23442, 25221, 25754, 25766, 24867, 23667, 23126, 22766, 22831, 
    23090, 23543, 24547, 25518, 26889, 25289, 26887, 26940, 26404, 25962, 
    25196, 24487,
  24829, 24944, 26435, 26444, 25956, 24889, 23645, 23060, 22851, 22815, 
    22998, 23513, 24431, 25604, 26637, 26797, 27495, 26979, 26488, 25901, 
    25172, 24602,
  25978, 26068, 26645, 26568, 25943, 24837, 23622, 23118, 22875, 22853, 
    22954, 23556, 24542, 25713, 26993, 27010, 27416, 26899, 26346, 25824, 
    25123, 24650,
  26408, 26543, 26628, 26538, 25891, 24773, 23580, 23048, 22833, 22828, 
    23081, 23690, 24408, 25806, 26950, 26992, 27424, 26822, 26259, 25638, 
    25054, 24544,
  26238, 26417, 26598, 26490, 25891, 24719, 23539, 23068, 22837, 22882, 
    23055, 23680, 24531, 25868, 26910, 27007, 27406, 26809, 26260, 25740, 
    25054, 24458,
  25710, 25867, 26552, 26451, 25826, 24722, 23541, 23088, 22831, 22874, 
    23138, 23614, 24579, 25759, 26822, 26926, 27373, 26793, 26274, 25665, 
    25049, 24412,
  24974, 25086, 26463, 26356, 25807, 24646, 23496, 23053, 22882, 22869, 
    23083, 23628, 24608, 25793, 26793, 26862, 27300, 26769, 26269, 25665, 
    24998, 24435,
  24132, 24227, 26100, 26206, 25668, 24622, 23470, 23031, 22887, 22879, 
    23087, 23565, 24519, 25819, 26881, 26531, 27332, 26769, 26295, 25672, 
    24940, 24429,
  23254, 23418, 25401, 25781, 25501, 24510, 23442, 23059, 22868, 22869, 
    23173, 23590, 24578, 25743, 27247, 25622, 27085, 26718, 26285, 25732, 
    24979, 24389,
  22445, 22724, 24774, 25430, 25394, 24458, 23405, 23076, 22893, 22948, 
    23023, 23674, 24642, 25739, 26928, 24410, 26440, 26646, 26188, 25694, 
    24987, 24383,
  21772, 22106, 24606, 25306, 25336, 24380, 23401, 22971, 22864, 22882, 
    23191, 23675, 24733, 25992, 27279, 23744, 26258, 26570, 26197, 25706, 
    25083, 24437,
  21154, 21439, 24649, 25371, 25243, 24332, 23349, 22985, 22869, 22927, 
    23098, 23618, 24754, 25863, 26771, 23556, 26316, 26597, 26219, 25776, 
    25122, 24464,
  20377, 20551, 24669, 25377, 25274, 24267, 23309, 22951, 22907, 22962, 
    23197, 23714, 24670, 26077, 26775, 23357, 26250, 26574, 26223, 25723, 
    25150, 24592,
  19394, 19468, 24643, 25380, 25212, 24246, 23267, 22968, 22866, 22959, 
    23310, 23701, 24790, 25926, 27232, 23269, 26357, 26561, 26151, 25604, 
    25062, 24554,
  18559, 18500, 24518, 25328, 25147, 24220, 23233, 22972, 22861, 23003, 
    23265, 23753, 24896, 25979, 26890, 23209, 26518, 26554, 26135, 25575, 
    24982, 24464,
  18373, 18053, 24610, 25350, 25132, 24182, 23177, 22912, 22932, 22918, 
    23213, 23824, 24707, 26262, 27212, 23070, 26704, 26422, 25943, 25465, 
    24737, 24012,
  18704, 18078, 24652, 25422, 25080, 24080, 23146, 22931, 22850, 22947, 
    23282, 23823, 24921, 26216, 26980, 22975, 26467, 26187, 25739, 25065, 
    24346, 23768,
  19393, 18543, 24747, 25197, 24886, 23841, 22998, 22769, 22794, 22950, 
    23280, 23855, 24828, 26270, 27159, 22676, 25269, 24949, 24708, 24351, 
    23790, 23345,
  28037, 28050, 27861, 27181, 25842, 24149, 22739, 22274, 22136, 22527, 
    22954, 23570, 24787, 25910, 26772, 28544, 28871, 27982, 27434, 26883, 
    26023, 25189,
  28027, 28041, 27888, 27299, 25978, 24284, 22769, 22306, 22144, 22483, 
    22930, 23672, 24584, 25753, 26373, 28582, 28960, 28022, 27470, 26852, 
    26055, 25142,
  27996, 28027, 27932, 27313, 26067, 24399, 22828, 22323, 22151, 22594, 
    22853, 23625, 24525, 25842, 26760, 28455, 28828, 27946, 27347, 26703, 
    25942, 25095,
  27915, 27983, 27719, 27306, 26148, 24517, 22929, 22371, 22157, 22423, 
    22862, 23467, 24507, 25887, 26478, 28236, 28680, 27857, 27288, 26783, 
    25910, 25007,
  27874, 27966, 27701, 27307, 26267, 24580, 23028, 22410, 22201, 22428, 
    22874, 23542, 24587, 25673, 26452, 28108, 28567, 27869, 27193, 26590, 
    25790, 24813,
  27860, 27965, 27650, 27340, 26265, 24689, 23075, 22422, 22201, 22489, 
    22767, 23492, 24460, 25707, 26607, 28096, 28503, 27857, 27221, 26572, 
    25732, 24860,
  27885, 27982, 27701, 27400, 26386, 24732, 23132, 22449, 22200, 22400, 
    22779, 23472, 24501, 25844, 26532, 28194, 28635, 27853, 27260, 26528, 
    25676, 24700,
  27956, 28045, 27860, 27501, 26490, 24868, 23216, 22526, 22223, 22516, 
    22901, 23435, 24408, 25793, 26315, 28350, 28851, 27881, 27183, 26503, 
    25574, 24431,
  28033, 28133, 27871, 27559, 26567, 24917, 23275, 22578, 22184, 22458, 
    22825, 23482, 24436, 25589, 26250, 28458, 28863, 27869, 27111, 26329, 
    25428, 24518,
  28053, 28187, 27943, 27617, 26616, 24992, 23311, 22569, 22242, 22438, 
    22776, 23482, 24334, 25737, 26483, 28394, 28796, 27735, 26971, 26194, 
    25237, 24299,
  28008, 28169, 27784, 27518, 26634, 25000, 23365, 22556, 22248, 22397, 
    22837, 23408, 24399, 25591, 26574, 28310, 28709, 27678, 26783, 26019, 
    25019, 24050,
  27936, 28106, 27685, 27422, 26591, 25073, 23407, 22601, 22243, 22468, 
    22800, 23434, 24363, 25709, 26557, 28121, 28482, 27530, 26712, 25872, 
    24865, 24028,
  27852, 28015, 27584, 27369, 26628, 25113, 23420, 22678, 22249, 22419, 
    22751, 23382, 24264, 25519, 26439, 28013, 28462, 27618, 26840, 25869, 
    24920, 24141,
  27759, 27897, 27576, 27386, 26682, 25197, 23534, 22703, 22300, 22461, 
    22798, 23348, 24340, 25462, 26432, 28020, 28583, 27765, 26953, 26054, 
    24969, 24172,
  27649, 27778, 27579, 27339, 26650, 25251, 23536, 22729, 22256, 22510, 
    22822, 23347, 24257, 25467, 26647, 27916, 28488, 27721, 26894, 25964, 
    25010, 24181,
  27554, 27693, 27407, 27285, 26674, 25259, 23601, 22760, 22297, 22462, 
    22795, 23479, 24313, 25418, 26997, 27723, 28231, 27560, 26754, 25924, 
    25053, 24199,
  27505, 27667, 27198, 27151, 26570, 25209, 23601, 22740, 22284, 22446, 
    22754, 23376, 24279, 25456, 26737, 27550, 28013, 27316, 26541, 25768, 
    24949, 24231,
  27521, 27688, 27271, 27175, 26657, 25324, 23703, 22821, 22339, 22418, 
    22822, 23413, 24285, 25362, 26413, 27586, 28019, 27263, 26382, 25612, 
    24910, 24255,
  27574, 27732, 27422, 27363, 26712, 25412, 23722, 22839, 22365, 22455, 
    22824, 23367, 24388, 25604, 26673, 27839, 28140, 27112, 26341, 25642, 
    24959, 24267,
  27633, 27781, 27546, 27378, 26795, 25429, 23761, 22912, 22364, 22422, 
    22819, 23470, 24343, 25399, 26376, 27962, 28144, 26926, 26126, 25510, 
    24865, 24255,
  27662, 27828, 27553, 27366, 26806, 25462, 23806, 22910, 22393, 22452, 
    22934, 23370, 24247, 25535, 26618, 27974, 28090, 26824, 26094, 25400, 
    24699, 24141,
  27670, 27861, 27516, 27372, 26739, 25476, 23795, 22915, 22400, 22448, 
    22818, 23253, 24192, 25671, 26191, 27900, 27987, 26757, 26059, 25438, 
    24762, 24026,
  27668, 27856, 27399, 27226, 26707, 25435, 23847, 22954, 22434, 22437, 
    22764, 23375, 24228, 25565, 26493, 27784, 27785, 26759, 26054, 25455, 
    24743, 24104,
  27624, 27775, 27291, 27156, 26661, 25443, 23860, 22963, 22417, 22501, 
    22790, 23399, 24226, 25307, 26863, 27668, 27575, 26632, 26015, 25448, 
    24773, 24191,
  27484, 27554, 27273, 27214, 26641, 25438, 23895, 23001, 22422, 22437, 
    22824, 23357, 24152, 25338, 26448, 27709, 27599, 26629, 25965, 25440, 
    24746, 24054,
  27220, 27196, 27275, 27188, 26701, 25493, 23896, 23004, 22462, 22425, 
    22750, 23320, 24201, 25403, 26310, 27694, 27640, 26597, 25999, 25377, 
    24724, 24080,
  26889, 26790, 26986, 27007, 26601, 25448, 23886, 23035, 22498, 22471, 
    22737, 23415, 24128, 25275, 26289, 27444, 27598, 26569, 25947, 25381, 
    24774, 24105,
  26611, 26490, 26660, 26813, 26541, 25473, 23924, 23010, 22529, 22451, 
    22857, 23330, 24170, 25490, 26478, 27104, 27379, 26525, 25924, 25366, 
    24766, 24078,
  26494, 26382, 26550, 26772, 26482, 25454, 23978, 23056, 22506, 22459, 
    22782, 23369, 24243, 25267, 26646, 26971, 27300, 26447, 25906, 25371, 
    24727, 24098,
  26562, 26465, 26701, 26846, 26541, 25524, 23994, 23056, 22508, 22436, 
    22796, 23335, 24126, 25235, 26609, 27112, 27353, 26393, 25841, 25289, 
    24695, 24024,
  26733, 26655, 26904, 26958, 26592, 25556, 24054, 23127, 22560, 22487, 
    22714, 23268, 24315, 25142, 26281, 27310, 27365, 26440, 25872, 25231, 
    24707, 24066,
  26898, 26860, 26987, 26966, 26603, 25504, 23996, 23075, 22554, 22495, 
    22707, 23393, 24241, 25127, 26311, 27316, 27333, 26407, 25829, 25244, 
    24695, 24133,
  26991, 26994, 26843, 26897, 26605, 25540, 24004, 23112, 22547, 22481, 
    22831, 23420, 24170, 25364, 26525, 27208, 27191, 26325, 25781, 25206, 
    24638, 24012,
  27026, 27034, 26837, 26916, 26563, 25521, 24063, 23112, 22564, 22488, 
    22783, 23350, 24161, 25317, 26563, 27222, 27160, 26266, 25744, 25275, 
    24682, 24039,
  27033, 27028, 26924, 26956, 26609, 25559, 24024, 23118, 22594, 22479, 
    22789, 23379, 24172, 25404, 26464, 27329, 27062, 26197, 25725, 25232, 
    24617, 24140,
  27019, 27019, 26994, 27000, 26603, 25524, 24056, 23201, 22581, 22479, 
    22755, 23341, 24093, 25272, 26157, 27397, 27015, 26175, 25676, 25171, 
    24553, 24098,
  26979, 27015, 26976, 26970, 26516, 25529, 24062, 23217, 22615, 22479, 
    22826, 23280, 24243, 25325, 26479, 27329, 26820, 26131, 25682, 25158, 
    24604, 24094,
  26919, 26983, 26894, 26839, 26507, 25523, 24069, 23200, 22594, 22568, 
    22745, 23272, 24097, 25265, 26769, 27112, 26650, 26144, 25676, 25238, 
    24623, 24054,
  26839, 26916, 26781, 26743, 26399, 25450, 24087, 23142, 22612, 22464, 
    22771, 23286, 24162, 25512, 26416, 26815, 26407, 26001, 25648, 25219, 
    24649, 23995,
  26742, 26816, 26593, 26518, 26276, 25404, 24020, 23169, 22641, 22468, 
    22750, 23258, 24083, 25323, 26475, 26471, 25916, 25788, 25524, 25237, 
    24624, 24071,
  26618, 26689, 26481, 26401, 26204, 25347, 24040, 23221, 22591, 22477, 
    22768, 23234, 24189, 25211, 26097, 26306, 25684, 25779, 25585, 25131, 
    24567, 23978,
  26478, 26541, 26369, 26424, 26094, 25329, 24059, 23198, 22672, 22482, 
    22814, 23320, 24154, 25289, 26157, 26239, 25993, 25966, 25694, 25249, 
    24741, 24020,
  26350, 26407, 26259, 26354, 26110, 25343, 24048, 23199, 22667, 22583, 
    22824, 23296, 24149, 25051, 26301, 26193, 26119, 25999, 25715, 25152, 
    24588, 24121,
  26590, 26507, 26641, 26515, 26247, 25304, 24034, 23131, 22598, 22536, 
    22787, 23221, 24013, 25260, 26335, 26401, 25664, 25787, 25565, 25168, 
    24620, 24082,
  26301, 26359, 26371, 26416, 26218, 25328, 24095, 23243, 22642, 22537, 
    22751, 23282, 24188, 25321, 26588, 26200, 25849, 25923, 25688, 25176, 
    24658, 24093,
  26408, 26471, 26469, 26507, 26228, 25399, 24067, 23230, 22663, 22526, 
    22865, 23299, 24250, 25296, 26424, 26338, 26093, 26001, 25713, 25308, 
    24722, 24108,
  26542, 26602, 26615, 26612, 26304, 25454, 24065, 23223, 22684, 22517, 
    22740, 23375, 24109, 25412, 26265, 26496, 25993, 25928, 25621, 25279, 
    24677, 24058,
  26647, 26697, 26644, 26653, 26300, 25426, 24076, 23208, 22682, 22544, 
    22837, 23294, 24248, 25443, 26309, 26516, 25982, 25959, 25644, 25274, 
    24707, 24137,
  26694, 26750, 26634, 26624, 26304, 25387, 24062, 23275, 22722, 22495, 
    22764, 23276, 24032, 25402, 26497, 26504, 26228, 26144, 25772, 25345, 
    24809, 24176,
  26705, 26777, 26565, 26575, 26286, 25388, 24045, 23261, 22672, 22500, 
    22744, 23276, 24225, 25253, 26408, 26403, 26182, 26041, 25770, 25281, 
    24688, 24189,
  26982, 26934, 26826, 26743, 26287, 25352, 24030, 23181, 22636, 22550, 
    22815, 23310, 24027, 25337, 26507, 26457, 25714, 25607, 25454, 25156, 
    24665, 24122,
  26950, 26902, 26938, 26749, 26342, 25405, 24044, 23163, 22616, 22561, 
    22767, 23282, 24245, 25321, 26324, 26557, 25645, 25685, 25461, 25112, 
    24633, 24109,
  26561, 26649, 26675, 26654, 26300, 25429, 24091, 23224, 22718, 22651, 
    22840, 23312, 24079, 25167, 26641, 26595, 26159, 25851, 25594, 25220, 
    24662, 24123,
  26366, 26452, 26585, 26640, 26318, 25386, 24058, 23243, 22727, 22604, 
    22899, 23269, 24155, 25426, 26585, 26676, 26118, 25774, 25540, 25191, 
    24560, 24001,
  26048, 26133, 26450, 26476, 26270, 25370, 24024, 23270, 22719, 22580, 
    22870, 23278, 24280, 25382, 26438, 26453, 25931, 25731, 25486, 25184, 
    24566, 24050,
  25655, 25745, 26143, 26294, 26211, 25324, 24051, 23226, 22754, 22581, 
    22889, 23296, 24159, 25385, 26550, 26141, 25558, 25562, 25407, 25122, 
    24605, 24002,
  25324, 25429, 25917, 26147, 26150, 25377, 24042, 23233, 22695, 22619, 
    22863, 23342, 24171, 25311, 26344, 25934, 26049, 25863, 25599, 25224, 
    24650, 24150,
  25233, 25346, 25744, 26116, 26124, 25310, 24032, 23197, 22684, 22620, 
    22921, 23306, 24312, 25289, 26193, 25904, 26406, 26085, 25675, 25218, 
    24739, 24017,
  25476, 25601, 26012, 26251, 26158, 25363, 23971, 23248, 22719, 22652, 
    22856, 23301, 24208, 25418, 26601, 26194, 26896, 26365, 25813, 25379, 
    24784, 24178,
  25988, 26130, 26513, 26625, 26393, 25432, 23997, 23225, 22767, 22698, 
    22815, 23425, 24335, 25219, 26494, 26791, 27313, 26578, 25984, 25424, 
    24671, 24138,
  26597, 26770, 27006, 26873, 26471, 25413, 23977, 23226, 22742, 22687, 
    22895, 23359, 24097, 25567, 26394, 27371, 27645, 26649, 25968, 25348, 
    24699, 24159,
  27097, 27320, 27237, 27068, 26546, 25448, 23998, 23232, 22762, 22652, 
    22843, 23321, 24171, 25490, 26450, 27588, 27723, 26732, 25990, 25350, 
    24636, 24174,
  27384, 27650, 27251, 27060, 26522, 25382, 23978, 23232, 22762, 22670, 
    22925, 23289, 24397, 25474, 26135, 27579, 27656, 26759, 26019, 25407, 
    24657, 24090,
  27483, 27751, 27173, 27024, 26513, 25386, 23971, 23207, 22762, 22658, 
    22925, 23344, 24346, 25423, 26525, 27538, 27742, 26829, 26164, 25407, 
    24682, 24132,
  27473, 27719, 27145, 27006, 26475, 25384, 23976, 23191, 22786, 22705, 
    22958, 23426, 24358, 25462, 26535, 27526, 27655, 26829, 26136, 25388, 
    24760, 24132,
  27423, 27651, 27194, 26922, 26468, 25349, 23924, 23184, 22754, 22756, 
    22882, 23394, 24155, 25378, 26488, 27536, 27747, 26915, 26160, 25425, 
    24728, 24153,
  27366, 27596, 27196, 26993, 26418, 25367, 23922, 23194, 22777, 22695, 
    22923, 23487, 24316, 25517, 26561, 27500, 27846, 26914, 26178, 25474, 
    24729, 24113,
  27296, 27553, 27101, 26969, 26438, 25351, 23912, 23177, 22770, 22754, 
    22852, 23379, 24199, 25395, 26215, 27419, 27838, 26975, 26206, 25532, 
    24755, 24190,
  27215, 27495, 26997, 26845, 26366, 25265, 23909, 23175, 22756, 22724, 
    22855, 23293, 24357, 25625, 26768, 27246, 27618, 27012, 26308, 25517, 
    24750, 24204,
  27142, 27394, 26867, 26781, 26308, 25242, 23886, 23177, 22770, 22701, 
    23052, 23385, 24340, 25324, 26757, 27159, 27505, 26994, 26339, 25558, 
    24834, 24239,
  27023, 27202, 26766, 26711, 26271, 25165, 23846, 23131, 22792, 22734, 
    23015, 23401, 24265, 25415, 26675, 27091, 27421, 26904, 26291, 25448, 
    24754, 24053,
  26689, 26788, 26756, 26684, 26195, 25120, 23798, 23148, 22778, 22731, 
    22967, 23337, 24303, 25427, 26536, 27016, 27400, 26889, 26328, 25601, 
    24869, 24217,
  25873, 25943, 26662, 26619, 26189, 25108, 23824, 23178, 22788, 22723, 
    22897, 23422, 24426, 25446, 26816, 27047, 27466, 26966, 26361, 25732, 
    24846, 24206,
  24438, 24536, 26116, 26325, 25999, 25070, 23786, 23139, 22798, 22742, 
    23016, 23440, 24380, 25890, 26682, 26734, 27501, 26999, 26422, 25793, 
    24975, 24273,
  22600, 22785, 24749, 25456, 25707, 24957, 23723, 23135, 22768, 22789, 
    22956, 23542, 24298, 25504, 26474, 25312, 27089, 27040, 26457, 25789, 
    25060, 24287,
  21011, 21290, 22942, 24487, 25324, 24826, 23701, 23101, 22807, 22782, 
    23031, 23497, 24256, 25651, 26667, 23012, 25626, 26808, 26436, 25907, 
    25129, 24417,
  20393, 20735, 22122, 24049, 25171, 24817, 23701, 23096, 22793, 22727, 
    22954, 23529, 24473, 25579, 26778, 21570, 25037, 26754, 26415, 25941, 
    25220, 24423,
  21088, 21376, 23117, 24602, 25391, 24806, 23693, 23106, 22818, 22792, 
    22969, 23549, 24336, 25639, 26701, 22478, 25355, 26831, 26434, 25844, 
    25215, 24491,
  22709, 22865, 25194, 25706, 25724, 24868, 23662, 23087, 22895, 22787, 
    23043, 23511, 24464, 25529, 26829, 25137, 26953, 26943, 26429, 25840, 
    25224, 24659,
  24449, 24467, 26414, 26439, 25956, 24865, 23663, 23086, 22848, 22800, 
    23065, 23576, 24357, 25676, 26718, 26807, 27535, 26946, 26451, 25959, 
    25333, 24674,
  25556, 25570, 26654, 26525, 25950, 24838, 23629, 23100, 22893, 22823, 
    23055, 23506, 24651, 25768, 26724, 27026, 27406, 26909, 26392, 25837, 
    25208, 24649,
  25813, 25898, 26560, 26484, 25835, 24752, 23563, 23069, 22854, 22856, 
    23031, 23526, 24525, 25576, 26550, 26983, 27378, 26925, 26394, 25902, 
    25273, 24683,
  25417, 25568, 26424, 26409, 25819, 24672, 23565, 23100, 22847, 22849, 
    23128, 23506, 24468, 25769, 26672, 26909, 27298, 26885, 26354, 25822, 
    25172, 24645,
  24699, 24847, 26313, 26312, 25753, 24650, 23524, 23040, 22858, 22861, 
    23069, 23569, 24428, 25788, 26662, 26775, 27283, 26825, 26347, 25834, 
    25076, 24599,
  23866, 23998, 26126, 26136, 25716, 24571, 23512, 23041, 22856, 22899, 
    23078, 23567, 24646, 25784, 26601, 26571, 27265, 26728, 26313, 25772, 
    25076, 24326,
  23049, 23194, 25443, 25826, 25562, 24545, 23426, 23054, 22885, 22884, 
    23043, 23649, 24631, 25906, 26729, 25865, 27072, 26721, 26250, 25791, 
    25076, 24428,
  22327, 22553, 24584, 25405, 25405, 24477, 23433, 23044, 22874, 22877, 
    23030, 23657, 24728, 25747, 26557, 24500, 26503, 26678, 26213, 25708, 
    25076, 24388,
  21792, 22108, 24396, 25178, 25339, 24425, 23382, 23031, 22887, 22895, 
    23110, 23626, 24666, 25951, 26778, 23554, 25982, 26656, 26234, 25751, 
    25085, 24522,
  21454, 21778, 24626, 25336, 25317, 24339, 23404, 22988, 22882, 22870, 
    23110, 23650, 24616, 25911, 26815, 23579, 26248, 26653, 26262, 25888, 
    25060, 24489,
  21145, 21383, 24747, 25419, 25268, 24331, 23364, 22976, 22893, 22895, 
    23106, 23712, 24541, 25950, 27029, 23639, 26244, 26700, 26285, 25963, 
    25233, 24703,
  20583, 20703, 24778, 25420, 25275, 24254, 23307, 22967, 22884, 22926, 
    23216, 23669, 24735, 26131, 27203, 23515, 26303, 26641, 26241, 25768, 
    25210, 24617,
  19687, 19737, 24756, 25429, 25197, 24233, 23258, 22962, 22834, 22906, 
    23181, 23732, 24759, 25966, 26828, 23426, 26447, 26636, 26196, 25648, 
    25129, 24667,
  18802, 18765, 24518, 25360, 25151, 24143, 23200, 22978, 22862, 22898, 
    23093, 23794, 24742, 26033, 26623, 23113, 26509, 26614, 26200, 25725, 
    25061, 24510,
  18454, 18183, 24539, 25332, 25133, 24114, 23186, 22926, 22908, 22886, 
    23226, 23731, 24733, 26228, 27015, 22729, 26547, 26512, 26097, 25505, 
    24842, 24272,
  18595, 18017, 24687, 25325, 25048, 24009, 23120, 22939, 22865, 22946, 
    23224, 23879, 24829, 26147, 27059, 22539, 26383, 26362, 25866, 25253, 
    24545, 23854,
  18758, 18014, 24820, 25366, 25057, 23940, 23104, 22896, 22859, 22953, 
    23268, 23777, 24987, 26099, 26723, 22493, 25870, 25653, 25212, 24732, 
    24176, 23602,
  28041, 28081, 27897, 27242, 25882, 24169, 22737, 22276, 22172, 22509, 
    22958, 23671, 24554, 25894, 26732, 28546, 28885, 28038, 27440, 26858, 
    26031, 25152,
  28029, 28073, 27932, 27322, 25956, 24271, 22789, 22270, 22137, 22493, 
    22859, 23601, 24684, 25782, 26750, 28529, 28919, 27941, 27413, 26846, 
    25974, 25052,
  27995, 28060, 27928, 27328, 26107, 24382, 22872, 22322, 22161, 22456, 
    22853, 23544, 24515, 25926, 26313, 28486, 28849, 27951, 27318, 26759, 
    25854, 24906,
  27914, 28013, 27815, 27321, 26159, 24501, 22972, 22355, 22179, 22485, 
    22837, 23599, 24549, 25815, 26856, 28278, 28657, 27826, 27225, 26641, 
    25816, 24892,
  27874, 27988, 27746, 27271, 26204, 24591, 22984, 22400, 22159, 22493, 
    22789, 23587, 24360, 25615, 26953, 28133, 28607, 27832, 27197, 26578, 
    25753, 24850,
  27853, 27973, 27675, 27307, 26281, 24676, 23090, 22450, 22194, 22457, 
    22784, 23581, 24393, 25801, 26309, 28054, 28480, 27913, 27199, 26603, 
    25753, 24790,
  27866, 27972, 27744, 27382, 26404, 24745, 23162, 22451, 22211, 22459, 
    22914, 23506, 24554, 25698, 26590, 28101, 28612, 27901, 27232, 26528, 
    25638, 24771,
  27924, 28021, 27881, 27468, 26453, 24852, 23221, 22510, 22260, 22451, 
    22868, 23493, 24323, 25636, 26588, 28232, 28759, 27915, 27175, 26459, 
    25588, 24608,
  27997, 28108, 27867, 27497, 26544, 24960, 23284, 22574, 22224, 22482, 
    22760, 23512, 24472, 25595, 26684, 28321, 28735, 27797, 27041, 26349, 
    25404, 24515,
  28018, 28169, 27848, 27555, 26601, 25037, 23323, 22586, 22243, 22517, 
    22831, 23437, 24464, 25514, 26800, 28322, 28797, 27734, 26969, 26144, 
    25169, 24155,
  27966, 28152, 27734, 27523, 26660, 25068, 23426, 22659, 22242, 22456, 
    22822, 23480, 24364, 25504, 26629, 28182, 28629, 27654, 26898, 26000, 
    25078, 24120,
  27879, 28080, 27714, 27449, 26660, 25065, 23457, 22651, 22272, 22479, 
    22821, 23457, 24407, 25715, 26462, 28070, 28651, 27730, 26924, 26151, 
    25096, 24112,
  27782, 27985, 27606, 27474, 26659, 25122, 23525, 22721, 22295, 22453, 
    22832, 23518, 24378, 25557, 26623, 28028, 28533, 27775, 27051, 26185, 
    25176, 24325,
  27693, 27871, 27568, 27401, 26657, 25214, 23539, 22714, 22325, 22457, 
    22810, 23409, 24409, 25491, 26978, 28006, 28579, 27785, 27110, 26276, 
    25257, 24356,
  27604, 27761, 27499, 27350, 26609, 25253, 23543, 22773, 22261, 22445, 
    22794, 23385, 24284, 25435, 26628, 27872, 28403, 27632, 26879, 26033, 
    25107, 24325,
  27534, 27683, 27354, 27259, 26631, 25259, 23619, 22798, 22331, 22451, 
    22781, 23383, 24260, 25414, 26949, 27683, 28178, 27326, 26504, 25750, 
    24966, 24276,
  27504, 27664, 27315, 27210, 26604, 25304, 23613, 22837, 22403, 22456, 
    22868, 23337, 24325, 25503, 26658, 27546, 27990, 27134, 26347, 25654, 
    24982, 24462,
  27536, 27693, 27328, 27219, 26643, 25353, 23711, 22820, 22343, 22511, 
    22794, 23479, 24252, 25474, 26616, 27607, 27940, 26966, 26276, 25637, 
    24937, 24326,
  27599, 27739, 27507, 27369, 26747, 25395, 23703, 22861, 22346, 22485, 
    22791, 23430, 24159, 25225, 26221, 27895, 28148, 26951, 26263, 25548, 
    24936, 24243,
  27657, 27774, 27649, 27485, 26826, 25441, 23800, 22917, 22395, 22518, 
    22794, 23387, 24362, 25505, 26550, 28015, 28153, 26779, 26056, 25516, 
    24859, 24252,
  27671, 27795, 27556, 27382, 26800, 25412, 23791, 22923, 22386, 22529, 
    22747, 23405, 24263, 25454, 26616, 27921, 27999, 26736, 26072, 25381, 
    24821, 24224,
  27650, 27795, 27372, 27266, 26699, 25407, 23818, 22917, 22469, 22484, 
    22770, 23411, 24285, 25623, 26569, 27735, 27665, 26591, 25968, 25412, 
    24764, 24131,
  27607, 27756, 27306, 27151, 26661, 25397, 23849, 22981, 22429, 22461, 
    22799, 23345, 24343, 25371, 26708, 27566, 27488, 26512, 25935, 25380, 
    24743, 24136,
  27525, 27649, 27254, 27145, 26635, 25410, 23847, 22986, 22459, 22471, 
    22832, 23313, 24268, 25339, 26475, 27515, 27403, 26522, 25944, 25390, 
    24743, 24135,
  27368, 27423, 27287, 27200, 26663, 25452, 23907, 23036, 22468, 22517, 
    22753, 23350, 24184, 25511, 26603, 27588, 27395, 26556, 25976, 25397, 
    24779, 24065,
  27128, 27090, 27144, 27153, 26694, 25509, 23884, 23003, 22506, 22487, 
    22867, 23355, 24230, 25558, 26240, 27548, 27455, 26487, 25900, 25339, 
    24713, 24083,
  26854, 26738, 26827, 26957, 26644, 25479, 23912, 23075, 22482, 22475, 
    22787, 23428, 24229, 25243, 26425, 27240, 27245, 26400, 25835, 25318, 
    24718, 24082,
  26632, 26497, 26481, 26745, 26524, 25471, 23953, 23076, 22517, 22515, 
    22889, 23340, 24214, 25430, 26665, 26928, 27220, 26414, 25832, 25316, 
    24698, 24035,
  26534, 26427, 26529, 26794, 26546, 25513, 23951, 23099, 22523, 22483, 
    22791, 23314, 24154, 25203, 26484, 26865, 27066, 26228, 25808, 25265, 
    24658, 24081,
  26568, 26495, 26790, 26896, 26581, 25553, 23985, 23096, 22498, 22538, 
    22814, 23264, 24223, 25332, 26454, 27043, 26882, 26153, 25626, 25252, 
    24632, 23947,
  26666, 26610, 26978, 26968, 26606, 25565, 23972, 23102, 22577, 22512, 
    22814, 23371, 24183, 25346, 26368, 27151, 26694, 25947, 25560, 25162, 
    24601, 24143,
  26745, 26701, 26969, 26957, 26606, 25525, 23987, 23113, 22551, 22552, 
    22813, 23320, 24212, 25298, 26248, 27104, 26526, 25885, 25497, 25082, 
    24563, 24022,
  26761, 26725, 26808, 26850, 26576, 25513, 24048, 23147, 22614, 22514, 
    22801, 23442, 24207, 25504, 26559, 26954, 26415, 25775, 25455, 25087, 
    24595, 23969,
  26740, 26694, 26690, 26797, 26515, 25496, 24030, 23180, 22630, 22453, 
    22809, 23360, 24112, 25301, 26176, 26898, 26410, 25831, 25468, 25051, 
    24506, 23835,
  26711, 26660, 26689, 26797, 26498, 25526, 24036, 23194, 22614, 22532, 
    22777, 23324, 24261, 25323, 26338, 26903, 26454, 25906, 25578, 25158, 
    24606, 24023,
  26683, 26650, 26598, 26679, 26492, 25536, 24044, 23203, 22612, 22558, 
    22796, 23315, 24331, 25246, 26326, 26828, 26506, 26065, 25640, 25215, 
    24619, 23995,
  26646, 26653, 26675, 26682, 26444, 25465, 24056, 23187, 22629, 22547, 
    22785, 23308, 24132, 25456, 26681, 26774, 26473, 26064, 25668, 25238, 
    24644, 24138,
  26594, 26626, 26613, 26685, 26387, 25471, 24067, 23185, 22634, 22555, 
    22815, 23277, 24148, 25512, 26359, 26729, 26528, 26185, 25750, 25238, 
    24676, 24017,
  26512, 26553, 26629, 26614, 26350, 25434, 24050, 23206, 22652, 22512, 
    22800, 23294, 24174, 25324, 26447, 26558, 26335, 26124, 25694, 25168, 
    24606, 24093,
  26709, 26609, 26870, 26710, 26301, 25364, 24042, 23145, 22580, 22586, 
    22748, 23353, 24163, 25270, 26457, 26482, 25728, 25857, 25536, 25143, 
    24539, 24153,
  26530, 26429, 26698, 26538, 26204, 25358, 24018, 23121, 22597, 22469, 
    22819, 23262, 24022, 25198, 26207, 26301, 25603, 25707, 25474, 25081, 
    24571, 24146,
  26012, 26050, 26190, 26275, 26097, 25314, 24095, 23250, 22659, 22490, 
    22821, 23229, 24264, 25535, 26309, 26058, 25788, 25907, 25672, 25224, 
    24697, 24157,
  25842, 25889, 26143, 26251, 26136, 25389, 24059, 23272, 22707, 22541, 
    22850, 23311, 24237, 25336, 26415, 26019, 25884, 25982, 25631, 25158, 
    24717, 24084,
  26066, 25985, 26388, 26403, 26179, 25383, 24049, 23177, 22644, 22609, 
    22753, 23254, 24165, 25450, 26167, 26145, 25578, 25670, 25480, 25162, 
    24603, 24079,
  26091, 26015, 26396, 26422, 26164, 25372, 24053, 23156, 22626, 22503, 
    22727, 23416, 24187, 25098, 26260, 26117, 25329, 25641, 25459, 25149, 
    24654, 24079,
  26212, 26135, 26589, 26557, 26242, 25369, 24042, 23147, 22632, 22554, 
    22770, 23259, 24178, 25214, 26312, 26268, 25815, 25713, 25563, 25162, 
    24629, 24092,
  26377, 26290, 26731, 26646, 26299, 25420, 24074, 23183, 22632, 22549, 
    22824, 23294, 24039, 25247, 26151, 26321, 25771, 25678, 25522, 25187, 
    24603, 24099,
  26528, 26430, 26785, 26743, 26273, 25412, 24042, 23212, 22652, 22574, 
    22858, 23320, 24316, 25268, 26260, 26396, 25715, 25735, 25556, 25149, 
    24609, 24139,
  26348, 26377, 26501, 26550, 26256, 25401, 24117, 23268, 22706, 22634, 
    22849, 23393, 24086, 25389, 26362, 26240, 25831, 25876, 25618, 25307, 
    24709, 24233,
  26687, 26580, 26804, 26694, 26307, 25403, 24035, 23203, 22638, 22571, 
    22853, 23305, 24128, 25163, 26454, 26401, 25435, 25446, 25273, 25037, 
    24565, 24058,
  26681, 26577, 26817, 26756, 26293, 25392, 24025, 23171, 22685, 22569, 
    22864, 23335, 24225, 25329, 26072, 26399, 24794, 24926, 25011, 24863, 
    24469, 24099,
  26599, 26515, 26832, 26692, 26256, 25414, 24039, 23168, 22682, 22606, 
    22844, 23343, 23992, 25121, 26373, 26415, 24794, 24984, 25059, 24944, 
    24450, 23945,
  26426, 26377, 26746, 26700, 26287, 25395, 24025, 23198, 22647, 22589, 
    22787, 23315, 24126, 25296, 26520, 26499, 25086, 25100, 25135, 24913, 
    24545, 24065,
  25862, 25977, 26262, 26427, 26218, 25432, 24057, 23295, 22729, 22597, 
    22911, 23292, 24211, 25217, 26312, 26202, 25260, 25217, 25223, 25003, 
    24536, 24079,
  25795, 25772, 26388, 26476, 26224, 25344, 24049, 23183, 22723, 22626, 
    22804, 23267, 24163, 25314, 26378, 26215, 25124, 25013, 24983, 24826, 
    24361, 23905,
  25393, 25350, 26134, 26366, 26196, 25291, 24001, 23142, 22650, 22638, 
    22850, 23391, 24054, 25340, 26390, 25992, 25417, 25244, 25149, 24926, 
    24475, 24086,
  25074, 25014, 25929, 26225, 26165, 25291, 24046, 23169, 22706, 22666, 
    22916, 23445, 24035, 25513, 26240, 25757, 26082, 25764, 25446, 25112, 
    24476, 24119,
  24693, 24794, 25460, 25959, 26078, 25378, 24044, 23267, 22768, 22713, 
    22984, 23378, 24136, 25459, 26617, 25444, 26545, 26199, 25701, 25243, 
    24626, 24048,
  24973, 25101, 25693, 26065, 26112, 25403, 24043, 23236, 22739, 22670, 
    22847, 23440, 24269, 25379, 26534, 25718, 26816, 26478, 25943, 25372, 
    24793, 24168,
  25564, 25719, 26184, 26425, 26269, 25385, 23998, 23239, 22749, 22694, 
    23038, 23435, 24243, 25367, 26538, 26339, 27216, 26642, 25969, 25368, 
    24736, 24181,
  26294, 26471, 26865, 26813, 26447, 25425, 24017, 23270, 22796, 22640, 
    22852, 23343, 24215, 25337, 26350, 27118, 27566, 26697, 26022, 25385, 
    24726, 24115,
  26930, 27143, 27210, 27019, 26515, 25420, 23982, 23246, 22728, 22682, 
    22948, 23347, 24245, 25325, 26665, 27481, 27744, 26759, 26037, 25381, 
    24746, 24137,
  27329, 27592, 27226, 27004, 26496, 25385, 23959, 23179, 22737, 22706, 
    22911, 23443, 24209, 25442, 26518, 27537, 27713, 26880, 26135, 25481, 
    24798, 24195,
  27493, 27787, 27130, 27012, 26488, 25376, 24007, 23232, 22784, 22614, 
    22862, 23423, 24268, 25480, 26566, 27477, 27744, 26921, 26204, 25507, 
    24825, 24143,
  27506, 27810, 27146, 26993, 26460, 25393, 23963, 23216, 22756, 22701, 
    22962, 23395, 24091, 25600, 26677, 27432, 27725, 27037, 26197, 25581, 
    24774, 24229,
  27465, 27756, 27113, 27013, 26454, 25350, 23981, 23257, 22762, 22672, 
    22845, 23417, 24221, 25672, 26499, 27469, 27768, 27028, 26255, 25668, 
    24768, 24251,
  27412, 27675, 27087, 26968, 26429, 25390, 23934, 23208, 22785, 22743, 
    22898, 23352, 24365, 25417, 26542, 27406, 27753, 26992, 26300, 25685, 
    24915, 24250,
  27317, 27560, 27029, 26943, 26398, 25319, 23931, 23209, 22751, 22737, 
    23007, 23371, 24290, 25519, 26411, 27416, 27803, 27053, 26356, 25707, 
    24960, 24307,
  27147, 27378, 26940, 26820, 26366, 25302, 23928, 23198, 22837, 22774, 
    22953, 23552, 24329, 25455, 26485, 27313, 27725, 27062, 26279, 25610, 
    24892, 24281,
  26907, 27110, 26866, 26813, 26322, 25231, 23891, 23197, 22813, 22768, 
    22962, 23434, 24295, 25446, 26857, 27184, 27582, 26950, 26290, 25595, 
    24886, 24249,
  26569, 26735, 26795, 26724, 26286, 25239, 23854, 23165, 22826, 22773, 
    22967, 23460, 24393, 25518, 26701, 27123, 27535, 26976, 26263, 25778, 
    24934, 24317,
  26024, 26166, 26738, 26651, 26198, 25092, 23797, 23156, 22862, 22768, 
    23019, 23434, 24226, 25434, 26506, 27066, 27501, 26981, 26382, 25818, 
    25024, 24328,
  25067, 25237, 26435, 26469, 26115, 25078, 23801, 23115, 22779, 22770, 
    22983, 23442, 24305, 25586, 26274, 26908, 27375, 26913, 26373, 25782, 
    25058, 24357,
  23596, 23833, 25480, 25881, 25839, 25020, 23756, 23158, 22809, 22823, 
    23042, 23509, 24326, 25782, 26261, 26047, 27160, 26925, 26337, 25854, 
    25072, 24304,
  21829, 22150, 23701, 24812, 25514, 24885, 23773, 23160, 22840, 22762, 
    22962, 23484, 24352, 25525, 26782, 23990, 25902, 26807, 26413, 25919, 
    25207, 24479,
  20383, 20741, 22334, 24131, 25232, 24793, 23728, 23115, 22861, 22831, 
    22958, 23424, 24438, 25801, 26730, 22025, 25112, 26741, 26407, 25994, 
    25296, 24521,
  19921, 20253, 22142, 24019, 25190, 24826, 23703, 23131, 22818, 22809, 
    22991, 23501, 24434, 25600, 26641, 21366, 24964, 26724, 26449, 25929, 
    25349, 24667,
  20714, 20916, 23325, 24674, 25377, 24829, 23698, 23138, 22867, 22784, 
    23058, 23486, 24354, 25626, 26758, 22510, 25220, 26750, 26466, 25999, 
    25306, 24642,
  22324, 22364, 25243, 25829, 25787, 24849, 23662, 23134, 22827, 22754, 
    22945, 23496, 24311, 25719, 26740, 25215, 26954, 26949, 26462, 25932, 
    25302, 24623,
  23928, 23848, 26491, 26406, 25931, 24894, 23657, 23073, 22847, 22850, 
    23083, 23511, 24395, 25709, 26624, 26879, 27674, 27009, 26498, 25878, 
    25367, 24671,
  24801, 24753, 26515, 26438, 25947, 24831, 23590, 23061, 22863, 22888, 
    23076, 23503, 24468, 25468, 26930, 27013, 27451, 26943, 26473, 25899, 
    25318, 24706,
  24785, 24846, 26225, 26223, 25838, 24767, 23586, 23097, 22835, 22917, 
    23051, 23556, 24579, 25633, 26491, 26784, 27378, 26837, 26379, 25908, 
    25262, 24600,
  24160, 24322, 25885, 26019, 25725, 24698, 23535, 23090, 22858, 22877, 
    23120, 23564, 24606, 25799, 26919, 26529, 27331, 26788, 26325, 25784, 
    25140, 24595,
  23326, 23525, 25581, 25910, 25670, 24611, 23498, 23065, 22854, 22866, 
    23103, 23562, 24595, 25778, 26997, 26225, 27204, 26744, 26276, 25797, 
    25142, 24556,
  22524, 22745, 25284, 25661, 25510, 24594, 23475, 23082, 22829, 22840, 
    23025, 23610, 24589, 25703, 26953, 25734, 27074, 26712, 26187, 25741, 
    25034, 24343,
  21881, 22132, 24556, 25358, 25374, 24504, 23451, 23043, 22816, 22920, 
    23114, 23542, 24618, 25849, 26909, 24621, 26651, 26691, 26185, 25729, 
    25053, 24498,
  21453, 21756, 23928, 25027, 25287, 24494, 23452, 23031, 22885, 22953, 
    23085, 23639, 24665, 25838, 27316, 23317, 25866, 26597, 26254, 25727, 
    25073, 24445,
  21284, 21614, 24061, 25091, 25270, 24431, 23425, 23060, 22863, 22896, 
    23167, 23651, 24561, 25829, 26891, 23057, 26072, 26525, 26239, 25751, 
    25074, 24559,
  21314, 21594, 24591, 25317, 25297, 24322, 23360, 23023, 22866, 22949, 
    23185, 23698, 24727, 26172, 26932, 23640, 26207, 26600, 26247, 25825, 
    25183, 24446,
  21307, 21472, 24871, 25418, 25288, 24310, 23306, 23004, 22871, 22939, 
    23166, 23700, 24742, 25988, 26955, 23789, 26246, 26663, 26235, 25901, 
    25248, 24747,
  20939, 20994, 25006, 25463, 25258, 24285, 23278, 22995, 22857, 22951, 
    23214, 23715, 24683, 26023, 26551, 23793, 26329, 26640, 26205, 25780, 
    25193, 24501,
  20122, 20137, 24906, 25468, 25223, 24256, 23259, 22961, 22862, 22976, 
    23173, 23762, 24842, 26049, 27034, 23734, 26429, 26584, 26229, 25766, 
    25150, 24490,
  19196, 19155, 24673, 25387, 25145, 24116, 23215, 22959, 22895, 23003, 
    23228, 23825, 24628, 26020, 27114, 23171, 26535, 26548, 26165, 25688, 
    25151, 24580,
  18689, 18433, 24567, 25296, 25102, 24103, 23191, 22954, 22861, 22938, 
    23162, 23789, 24747, 26187, 27320, 22515, 26412, 26510, 26118, 25573, 
    24964, 24309,
  18633, 18075, 24671, 25386, 25059, 24071, 23110, 22979, 22854, 23048, 
    23176, 23740, 24824, 26382, 27192, 22360, 26323, 26475, 25954, 25370, 
    24718, 24018,
  18706, 17981, 24883, 25424, 25006, 23940, 23078, 22892, 22867, 22937, 
    23193, 23823, 24953, 26349, 27071, 22390, 26058, 25925, 25487, 24968, 
    24254, 23685,
  28066, 28084, 27919, 27266, 25882, 24171, 22712, 22278, 22221, 22528, 
    23004, 23627, 24740, 25947, 26587, 28563, 28903, 28069, 27519, 26899, 
    26055, 25089,
  28054, 28078, 27926, 27328, 26018, 24279, 22761, 22268, 22174, 22519, 
    22870, 23628, 24682, 25615, 26629, 28537, 28924, 28059, 27472, 26879, 
    26010, 25103,
  28020, 28071, 27868, 27432, 26101, 24410, 22899, 22348, 22178, 22478, 
    22898, 23493, 24666, 25956, 26585, 28558, 28841, 27961, 27369, 26756, 
    25916, 24903,
  27937, 28030, 27879, 27347, 26228, 24497, 22972, 22384, 22187, 22525, 
    22868, 23575, 24549, 25612, 26341, 28328, 28731, 27866, 27297, 26724, 
    25865, 25043,
  27891, 28011, 27747, 27295, 26273, 24593, 23012, 22373, 22181, 22522, 
    22850, 23580, 24555, 25755, 26387, 28211, 28593, 27834, 27207, 26662, 
    25789, 24761,
  27861, 27997, 27724, 27355, 26281, 24669, 23132, 22437, 22186, 22451, 
    22780, 23454, 24684, 25735, 26669, 28126, 28567, 27858, 27223, 26637, 
    25757, 24874,
  27860, 27987, 27659, 27369, 26403, 24790, 23148, 22473, 22213, 22518, 
    22947, 23558, 24468, 25830, 26741, 28126, 28579, 27860, 27297, 26600, 
    25701, 24734,
  27907, 28021, 27796, 27468, 26467, 24857, 23249, 22547, 22212, 22425, 
    22958, 23581, 24464, 25733, 26552, 28269, 28703, 27866, 27137, 26494, 
    25471, 24620,
  27975, 28092, 27835, 27518, 26513, 24957, 23274, 22508, 22249, 22442, 
    22829, 23401, 24226, 25641, 26590, 28296, 28790, 27799, 27030, 26257, 
    25364, 24453,
  27996, 28140, 27785, 27508, 26613, 24998, 23312, 22587, 22220, 22448, 
    22764, 23529, 24307, 25666, 26507, 28288, 28728, 27722, 26932, 26178, 
    25141, 24213,
  27937, 28109, 27791, 27479, 26637, 25087, 23371, 22619, 22252, 22430, 
    22854, 23458, 24257, 25545, 26594, 28254, 28703, 27765, 26874, 26121, 
    25133, 24265,
  27833, 28026, 27700, 27488, 26676, 25078, 23406, 22660, 22262, 22495, 
    22737, 23487, 24238, 25366, 26440, 28174, 28694, 27805, 27017, 26229, 
    25145, 24378,
  27723, 27933, 27563, 27426, 26650, 25178, 23525, 22700, 22320, 22492, 
    22820, 23415, 24402, 25751, 26457, 28050, 28557, 27741, 27000, 26250, 
    25155, 24390,
  27642, 27836, 27510, 27393, 26588, 25183, 23484, 22698, 22269, 22390, 
    22842, 23481, 24401, 25651, 26251, 27956, 28454, 27709, 26900, 26112, 
    25089, 24307,
  27578, 27745, 27447, 27307, 26647, 25201, 23576, 22742, 22286, 22407, 
    22801, 23373, 24208, 25435, 26607, 27825, 28153, 27368, 26572, 25849, 
    25010, 24236,
  27534, 27676, 27346, 27254, 26623, 25202, 23585, 22770, 22342, 22453, 
    22731, 23386, 24350, 25560, 26253, 27731, 28015, 27013, 26232, 25560, 
    24798, 24200,
  27516, 27655, 27271, 27247, 26624, 25281, 23662, 22862, 22370, 22490, 
    22761, 23416, 24274, 25321, 26596, 27675, 27914, 26826, 26150, 25503, 
    24828, 24218,
  27542, 27675, 27335, 27281, 26663, 25285, 23669, 22842, 22425, 22430, 
    22790, 23307, 24317, 25221, 26513, 27719, 27852, 26701, 26025, 25403, 
    24787, 24210,
  27587, 27707, 27478, 27343, 26675, 25332, 23717, 22845, 22384, 22402, 
    22769, 23386, 24193, 25484, 26451, 27898, 27935, 26651, 25976, 25451, 
    24883, 24235,
  27623, 27717, 27513, 27344, 26746, 25364, 23752, 22836, 22397, 22443, 
    22798, 23373, 24143, 25295, 26522, 27884, 27916, 26602, 25991, 25481, 
    24839, 24183,
  27620, 27707, 27370, 27195, 26711, 25418, 23801, 22949, 22412, 22479, 
    22808, 23336, 24343, 25562, 26445, 27778, 27755, 26508, 25888, 25390, 
    24812, 24162,
  27587, 27677, 27219, 27150, 26647, 25378, 23836, 22916, 22434, 22421, 
    22709, 23333, 24258, 25381, 26100, 27574, 27315, 26485, 25937, 25465, 
    24768, 24215,
  27529, 27616, 27211, 27082, 26615, 25368, 23832, 22962, 22467, 22415, 
    22840, 23359, 24274, 25295, 26477, 27480, 27306, 26428, 25959, 25414, 
    24825, 24134,
  27421, 27499, 27245, 27163, 26592, 25454, 23837, 22969, 22482, 22451, 
    22792, 23408, 24200, 25251, 26416, 27565, 27265, 26489, 25926, 25506, 
    24836, 24159,
  27251, 27290, 27195, 27151, 26621, 25454, 23859, 23000, 22429, 22508, 
    22765, 23348, 24371, 25446, 26443, 27591, 27438, 26500, 25897, 25382, 
    24687, 24062,
  27037, 27013, 26950, 26966, 26570, 25432, 23923, 23010, 22518, 22375, 
    22851, 23402, 24260, 25315, 26747, 27459, 27367, 26447, 25849, 25249, 
    24685, 23988,
  26834, 26746, 26689, 26829, 26519, 25489, 23920, 23039, 22496, 22458, 
    22834, 23269, 24165, 25241, 26544, 27087, 26976, 26179, 25728, 25353, 
    24626, 23993,
  26691, 26593, 26518, 26731, 26504, 25428, 23943, 23064, 22484, 22477, 
    22865, 23288, 24076, 25262, 26531, 26875, 26826, 26071, 25684, 25187, 
    24594, 23986,
  26638, 26579, 26579, 26766, 26500, 25501, 23969, 23089, 22524, 22483, 
    22778, 23386, 24129, 25219, 26133, 26929, 26778, 26029, 25535, 25169, 
    24523, 23872,
  26658, 26641, 26841, 26850, 26553, 25487, 23950, 23075, 22579, 22471, 
    22741, 23420, 24164, 25317, 26373, 27082, 26625, 25997, 25505, 25080, 
    24510, 23851,
  26694, 26688, 26906, 26906, 26552, 25463, 24007, 23063, 22573, 22468, 
    22728, 23303, 24140, 25362, 26734, 27087, 26281, 25669, 25378, 25053, 
    24496, 23974,
  26688, 26675, 26868, 26806, 26526, 25479, 23998, 23135, 22570, 22543, 
    22834, 23296, 24172, 25328, 26443, 26951, 25914, 25543, 25307, 25067, 
    24504, 23880,
  26624, 26602, 26627, 26722, 26462, 25479, 24002, 23128, 22610, 22499, 
    22773, 23319, 24197, 25306, 26116, 26834, 26083, 25654, 25417, 25034, 
    24516, 24033,
  26539, 26504, 26519, 26634, 26375, 25453, 24002, 23146, 22587, 22524, 
    22779, 23361, 24156, 25252, 26184, 26778, 26184, 25791, 25526, 25172, 
    24643, 24013,
  26469, 26436, 26461, 26632, 26391, 25427, 24036, 23134, 22574, 22468, 
    22807, 23271, 24117, 25504, 26682, 26700, 26278, 25881, 25526, 25191, 
    24521, 23940,
  26422, 26411, 26401, 26557, 26337, 25393, 24037, 23172, 22620, 22478, 
    22814, 23322, 24151, 25251, 26390, 26605, 26291, 25909, 25518, 25180, 
    24572, 23986,
  26383, 26406, 26354, 26484, 26341, 25434, 24050, 23180, 22645, 22504, 
    22779, 23322, 24194, 25503, 26213, 26545, 26316, 25937, 25587, 25247, 
    24585, 24009,
  26330, 26370, 26393, 26484, 26241, 25380, 24043, 23154, 22651, 22466, 
    22861, 23291, 23961, 25487, 26548, 26513, 26413, 26029, 25684, 25272, 
    24635, 24069,
  26224, 26274, 26326, 26446, 26197, 25363, 24047, 23182, 22633, 22528, 
    22813, 23254, 24199, 25399, 26213, 26377, 26171, 25938, 25629, 25290, 
    24674, 24144,
  26044, 26097, 26293, 26376, 26204, 25396, 24077, 23203, 22665, 22550, 
    22923, 23287, 24062, 25237, 26200, 26162, 25991, 25919, 25615, 25240, 
    24623, 24166,
  25796, 25848, 26138, 26287, 26116, 25367, 24062, 23186, 22659, 22538, 
    22793, 23251, 24147, 25162, 26396, 25979, 25809, 25846, 25621, 25146, 
    24643, 24060,
  25529, 25573, 26026, 26220, 26082, 25381, 24043, 23169, 22649, 22475, 
    22816, 23306, 24151, 25353, 26275, 26016, 25962, 25925, 25613, 25283, 
    24695, 24148,
  25307, 25354, 25924, 26193, 26121, 25355, 24025, 23229, 22697, 22564, 
    22828, 23270, 24119, 25330, 26197, 25935, 26075, 25978, 25660, 25241, 
    24664, 24110,
  25198, 25241, 25828, 26169, 26082, 25323, 24020, 23236, 22675, 22492, 
    22810, 23284, 24151, 25118, 26378, 25838, 25810, 25868, 25644, 25304, 
    24677, 24170,
  25526, 25421, 26138, 26241, 26113, 25304, 23997, 23128, 22634, 22482, 
    22743, 23189, 24087, 25324, 26135, 25984, 25483, 25695, 25539, 25140, 
    24524, 24110,
  25359, 25372, 25921, 26163, 26107, 25335, 24076, 23243, 22708, 22522, 
    22829, 23359, 24012, 25468, 26761, 25826, 25962, 25823, 25618, 25242, 
    24651, 24129,
  25547, 25555, 26087, 26224, 26129, 25297, 24109, 23204, 22749, 22581, 
    22839, 23336, 24050, 25185, 26270, 25897, 25904, 25821, 25601, 25232, 
    24695, 24187,
  26019, 25896, 26359, 26462, 26184, 25341, 24029, 23149, 22666, 22548, 
    22917, 23321, 24030, 25287, 26245, 26101, 25826, 25846, 25560, 25177, 
    24652, 24130,
  25884, 25891, 26041, 26269, 26153, 25339, 24034, 23275, 22705, 22617, 
    22814, 23323, 24296, 25312, 26357, 25995, 25991, 25972, 25663, 25335, 
    24674, 24111,
  25983, 25967, 26118, 26353, 26160, 25385, 24082, 23206, 22758, 22627, 
    22754, 23349, 24164, 25433, 26571, 26094, 25965, 25854, 25592, 25302, 
    24700, 24190,
  25983, 25957, 26306, 26398, 26233, 25386, 24057, 23252, 22708, 22607, 
    22820, 23351, 24083, 25301, 26393, 26133, 25574, 25487, 25443, 25230, 
    24655, 24223,
  26166, 26026, 26499, 26534, 26226, 25293, 24039, 23137, 22651, 22560, 
    22840, 23242, 24141, 25326, 26443, 26268, 25047, 25132, 25152, 24978, 
    24512, 24144,
  25935, 25845, 26316, 26416, 26154, 25304, 24018, 23137, 22654, 22623, 
    22734, 23298, 24084, 25410, 26165, 26101, 25010, 25081, 25118, 24978, 
    24614, 24097,
  25607, 25556, 26098, 26235, 26129, 25321, 24008, 23188, 22684, 22549, 
    22797, 23296, 24166, 25231, 26334, 25892, 25054, 25103, 25069, 24978, 
    24518, 24070,
  25213, 25164, 25951, 26190, 26144, 25299, 24005, 23140, 22637, 22632, 
    22783, 23362, 24084, 25291, 26325, 25782, 25209, 25262, 25145, 24997, 
    24461, 24030,
  24806, 24731, 25851, 26092, 26069, 25271, 23987, 23140, 22655, 22580, 
    22806, 23248, 24097, 25257, 26456, 25685, 25851, 25644, 25380, 25015, 
    24607, 23996,
  24490, 24396, 25707, 25988, 26026, 25282, 23997, 23161, 22681, 22594, 
    22883, 23263, 24109, 25138, 26326, 25546, 26279, 25970, 25553, 25190, 
    24601, 24084,
  24110, 24184, 25234, 25810, 25969, 25296, 24003, 23192, 22717, 22638, 
    22798, 23354, 24173, 25501, 26615, 25171, 26606, 26375, 25850, 25264, 
    24611, 24099,
  24404, 24522, 25337, 25857, 26000, 25309, 24001, 23223, 22759, 22687, 
    22897, 23276, 24260, 25345, 26101, 25253, 26666, 26510, 25910, 25301, 
    24740, 24092,
  25054, 25209, 25826, 26159, 26137, 25312, 24016, 23235, 22783, 22708, 
    22905, 23401, 24335, 25397, 26414, 25893, 26984, 26572, 25944, 25346, 
    24722, 24099,
  25900, 26073, 26594, 26654, 26325, 25340, 24017, 23230, 22737, 22665, 
    22857, 23387, 24144, 25305, 26225, 26895, 27522, 26765, 25991, 25400, 
    24673, 24160,
  26692, 26886, 27041, 26963, 26423, 25420, 23965, 23239, 22739, 22699, 
    22815, 23335, 24186, 25444, 26263, 27468, 27650, 26841, 26082, 25477, 
    24795, 24189,
  27242, 27478, 27190, 27010, 26456, 25429, 23970, 23246, 22807, 22649, 
    22870, 23426, 24253, 25335, 26525, 27495, 27762, 26890, 26153, 25422, 
    24764, 24193,
  27509, 27788, 27142, 26987, 26421, 25372, 23948, 23234, 22795, 22714, 
    22943, 23396, 24279, 25436, 26561, 27429, 27662, 27004, 26255, 25528, 
    24829, 24349,
  27561, 27867, 27094, 26984, 26478, 25381, 23905, 23253, 22784, 22660, 
    22911, 23425, 24259, 25547, 26685, 27479, 27674, 27069, 26290, 25577, 
    24893, 24301,
  27501, 27792, 27008, 26915, 26445, 25316, 23929, 23240, 22801, 22705, 
    22971, 23413, 24229, 25311, 26509, 27449, 27804, 27053, 26314, 25614, 
    24932, 24342,
  27381, 27613, 26957, 26916, 26431, 25287, 23921, 23212, 22834, 22728, 
    22982, 23424, 24277, 25457, 26339, 27334, 27666, 27031, 26310, 25669, 
    24939, 24301,
  27159, 27325, 26917, 26825, 26363, 25287, 23879, 23149, 22797, 22711, 
    23054, 23403, 24151, 25562, 26707, 27310, 27634, 27055, 26359, 25653, 
    24888, 24325,
  26778, 26911, 26937, 26822, 26265, 25248, 23886, 23167, 22775, 22728, 
    22940, 23520, 24253, 25388, 26413, 27249, 27581, 26934, 26323, 25631, 
    24941, 24259,
  26248, 26382, 26875, 26731, 26214, 25222, 23822, 23136, 22818, 22717, 
    23080, 23453, 24213, 25460, 26532, 27212, 27581, 26959, 26286, 25654, 
    24903, 24287,
  25611, 25775, 26603, 26585, 26140, 25129, 23815, 23173, 22801, 22870, 
    22943, 23451, 24302, 25381, 26691, 27060, 27565, 26957, 26315, 25681, 
    24964, 24349,
  24869, 25080, 26216, 26356, 26049, 25047, 23800, 23146, 22832, 22760, 
    22961, 23463, 24219, 25367, 26384, 26818, 27550, 26969, 26350, 25833, 
    25047, 24312,
  23906, 24188, 25838, 26149, 25969, 25049, 23812, 23197, 22766, 22770, 
    22990, 23510, 24424, 25347, 26608, 26521, 27410, 27004, 26452, 25847, 
    25145, 24469,
  22633, 22984, 24899, 25591, 25755, 24960, 23771, 23124, 22796, 22768, 
    22977, 23487, 24346, 25509, 26591, 25374, 26967, 26871, 26458, 25888, 
    25108, 24422,
  21187, 21585, 23491, 24764, 25431, 24865, 23756, 23168, 22859, 22818, 
    23035, 23429, 24323, 25570, 26584, 23277, 25482, 26753, 26451, 25997, 
    25339, 24611,
  20050, 20416, 22587, 24250, 25237, 24815, 23735, 23142, 22825, 22839, 
    22970, 23458, 24212, 25589, 26762, 21928, 25060, 26801, 26451, 25966, 
    25340, 24559,
  19754, 20021, 22458, 24179, 25223, 24834, 23711, 23105, 22838, 22806, 
    23075, 23469, 24306, 25649, 26718, 21619, 24943, 26697, 26369, 26006, 
    25297, 24545,
  20499, 20599, 23636, 24748, 25382, 24751, 23687, 23063, 22829, 22833, 
    23076, 23495, 24467, 25697, 26444, 22833, 25548, 26768, 26415, 25934, 
    25253, 24553,
  21865, 21822, 25445, 25845, 25810, 24828, 23660, 23112, 22850, 22817, 
    23109, 23591, 24304, 25860, 26496, 25437, 27146, 26959, 26438, 25929, 
    25300, 24674,
  23117, 23000, 26383, 26386, 25900, 24871, 23592, 23128, 22816, 22847, 
    23107, 23593, 24395, 25848, 26310, 26857, 27685, 26982, 26411, 25875, 
    25154, 24682,
  23633, 23589, 26104, 26187, 25794, 24771, 23562, 23104, 22847, 22841, 
    23009, 23598, 24511, 25751, 26604, 26731, 27401, 26824, 26380, 25921, 
    25214, 24717,
  23343, 23430, 25522, 25847, 25664, 24730, 23596, 23099, 22855, 22890, 
    23107, 23580, 24575, 25810, 26819, 26059, 27178, 26754, 26306, 25817, 
    25126, 24558,
  22584, 22791, 24845, 25503, 25492, 24661, 23553, 23097, 22848, 22871, 
    23113, 23596, 24584, 25743, 26922, 25350, 26850, 26697, 26273, 25775, 
    25114, 24519,
  21783, 22051, 24387, 25282, 25444, 24577, 23484, 23076, 22894, 22877, 
    23070, 23626, 24590, 25829, 27066, 24795, 26680, 26790, 26218, 25706, 
    25044, 24420,
  21173, 21478, 24082, 25092, 25350, 24551, 23451, 23072, 22880, 22889, 
    23183, 23652, 24501, 25791, 27088, 24147, 26357, 26657, 26232, 25706, 
    25051, 24428,
  20842, 21163, 23739, 24899, 25257, 24453, 23437, 23043, 22900, 22971, 
    23096, 23643, 24589, 25974, 26641, 23296, 25991, 26672, 26190, 25744, 
    25083, 24409,
  20793, 21116, 23628, 24840, 25233, 24424, 23390, 23045, 22901, 22904, 
    23094, 23688, 24648, 25831, 26676, 22575, 25726, 26585, 26195, 25717, 
    25064, 24363,
  21011, 21301, 24117, 25098, 25252, 24408, 23442, 23015, 22894, 22942, 
    23106, 23718, 24687, 25799, 26991, 22912, 26007, 26564, 26222, 25723, 
    24983, 24436,
  21377, 21586, 24734, 25380, 25331, 24369, 23401, 23045, 22868, 22934, 
    23189, 23708, 24567, 25960, 26841, 23692, 26248, 26683, 26257, 25791, 
    25193, 24557,
  21609, 21719, 25010, 25495, 25282, 24303, 23314, 22980, 22923, 22890, 
    23201, 23640, 24553, 25969, 26972, 23951, 26344, 26600, 26218, 25767, 
    25245, 24558,
  21381, 21420, 25117, 25561, 25226, 24274, 23292, 22993, 22911, 22893, 
    23138, 23665, 24838, 26055, 26847, 24056, 26334, 26585, 26140, 25814, 
    25120, 24504,
  20623, 20648, 25101, 25540, 25211, 24219, 23277, 22986, 22896, 22993, 
    23125, 23744, 24675, 25997, 27124, 24040, 26453, 26594, 26150, 25713, 
    25071, 24447,
  19667, 19643, 24743, 25396, 25127, 24148, 23195, 22934, 22871, 22917, 
    23140, 23828, 24779, 26136, 27013, 23313, 26553, 26566, 26085, 25653, 
    25054, 24377,
  19028, 18787, 24584, 25346, 25072, 24085, 23201, 22959, 22862, 22993, 
    23169, 23828, 24871, 26266, 26682, 22412, 26348, 26469, 26031, 25526, 
    24987, 24374,
  18796, 18249, 24810, 25396, 25050, 24028, 23159, 22958, 22904, 22927, 
    23254, 23769, 24910, 26096, 27232, 22485, 26377, 26435, 25985, 25404, 
    24735, 24056,
  18785, 18070, 25085, 25471, 24979, 23904, 23072, 22900, 22884, 22951, 
    23170, 23778, 24938, 26328, 26738, 22576, 26224, 26201, 25656, 25162, 
    24412, 23650,
  28095, 28087, 27906, 27239, 25891, 24183, 22679, 22282, 22178, 22432, 
    22914, 23654, 24674, 25814, 26480, 28581, 28925, 28045, 27515, 26965, 
    26013, 24974,
  28084, 28081, 27966, 27257, 25967, 24268, 22800, 22293, 22149, 22517, 
    22912, 23609, 24719, 25697, 26394, 28532, 28964, 28086, 27482, 26729, 
    25924, 24900,
  28050, 28074, 27945, 27312, 26092, 24396, 22810, 22263, 22137, 22465, 
    22906, 23570, 24628, 25840, 26604, 28559, 28944, 27973, 27428, 26772, 
    25894, 24867,
  27963, 28039, 27784, 27353, 26184, 24478, 22917, 22326, 22144, 22512, 
    22918, 23548, 24471, 25539, 26524, 28354, 28709, 27834, 27252, 26672, 
    25829, 24879,
  27910, 28030, 27694, 27295, 26230, 24600, 23023, 22394, 22156, 22472, 
    22962, 23594, 24482, 25834, 26457, 28211, 28596, 27774, 27156, 26499, 
    25671, 24658,
  27869, 28022, 27706, 27342, 26278, 24655, 23092, 22426, 22187, 22532, 
    22812, 23526, 24609, 25751, 26882, 28068, 28526, 27834, 27212, 26499, 
    25632, 24538,
  27854, 28005, 27712, 27337, 26354, 24699, 23124, 22427, 22196, 22518, 
    22926, 23504, 24475, 25597, 26507, 28119, 28563, 27881, 27191, 26425, 
    25596, 24632,
  27886, 28015, 27743, 27408, 26464, 24815, 23195, 22493, 22175, 22487, 
    22843, 23436, 24296, 25653, 26407, 28213, 28662, 27822, 27071, 26362, 
    25385, 24463,
  27943, 28058, 27840, 27479, 26510, 24912, 23229, 22547, 22179, 22421, 
    22847, 23421, 24428, 25662, 26725, 28299, 28762, 27803, 27040, 26244, 
    25246, 24290,
  27959, 28084, 27838, 27541, 26613, 24931, 23297, 22600, 22187, 22452, 
    22862, 23549, 24614, 25712, 26606, 28332, 28819, 27800, 27010, 26176, 
    25137, 24251,
  27898, 28039, 27801, 27522, 26581, 25023, 23410, 22626, 22247, 22406, 
    22751, 23501, 24257, 25612, 26497, 28285, 28794, 27806, 27001, 26243, 
    25206, 24203,
  27791, 27948, 27685, 27470, 26646, 25073, 23432, 22654, 22260, 22466, 
    22831, 23397, 24387, 25629, 26315, 28160, 28673, 27752, 26930, 26197, 
    25167, 24188,
  27683, 27858, 27594, 27368, 26630, 25158, 23450, 22704, 22301, 22460, 
    22783, 23415, 24328, 25577, 26256, 28041, 28515, 27603, 26885, 26038, 
    25082, 24133,
  27615, 27777, 27468, 27342, 26607, 25205, 23512, 22687, 22294, 22439, 
    22834, 23473, 24342, 25525, 26800, 27906, 28357, 27425, 26612, 25912, 
    25080, 24311,
  27574, 27707, 27381, 27276, 26600, 25171, 23546, 22740, 22343, 22429, 
    22855, 23395, 24372, 25295, 26249, 27806, 28018, 27128, 26326, 25661, 
    24803, 24147,
  27549, 27651, 27344, 27228, 26591, 25191, 23590, 22750, 22381, 22446, 
    22786, 23373, 24349, 25511, 26246, 27676, 27806, 26671, 25979, 25453, 
    24801, 24037,
  27529, 27631, 27276, 27190, 26529, 25220, 23635, 22779, 22353, 22440, 
    22824, 23425, 24207, 25661, 26448, 27547, 27232, 26284, 25773, 25333, 
    24678, 24217,
  27531, 27640, 27281, 27178, 26579, 25299, 23653, 22832, 22387, 22444, 
    22801, 23380, 24277, 25425, 26294, 27463, 27052, 26209, 25759, 25283, 
    24689, 24141,
  27540, 27651, 27384, 27225, 26632, 25307, 23680, 22884, 22379, 22444, 
    22775, 23271, 24309, 25394, 26760, 27578, 26860, 26260, 25779, 25375, 
    24783, 24153,
  27542, 27637, 27275, 27282, 26654, 25340, 23739, 22899, 22422, 22451, 
    22809, 23316, 24310, 25474, 26466, 27617, 27146, 26376, 25849, 25442, 
    24821, 24120,
  27523, 27605, 27264, 27225, 26625, 25392, 23809, 22899, 22400, 22467, 
    22797, 23406, 24406, 25519, 26512, 27581, 27335, 26433, 25891, 25351, 
    24751, 24127,
  27495, 27561, 27172, 27118, 26644, 25373, 23819, 22955, 22414, 22460, 
    22746, 23350, 24292, 25392, 26559, 27462, 27449, 26410, 25815, 25296, 
    24662, 24073,
  27443, 27491, 27183, 27123, 26609, 25359, 23826, 23025, 22476, 22434, 
    22790, 23452, 24192, 25371, 26457, 27516, 27382, 26426, 25914, 25332, 
    24707, 24118,
  27329, 27374, 27176, 27169, 26609, 25434, 23842, 22964, 22424, 22436, 
    22823, 23333, 24179, 25321, 26307, 27621, 27416, 26443, 25832, 25379, 
    24731, 24050,
  27155, 27192, 27048, 27041, 26580, 25426, 23901, 22986, 22503, 22415, 
    22749, 23332, 24280, 25401, 26583, 27555, 27496, 26404, 25825, 25362, 
    24582, 24074,
  26973, 26981, 26775, 26860, 26507, 25424, 23934, 22991, 22493, 22483, 
    22782, 23353, 24149, 25215, 26415, 27315, 27369, 26379, 25810, 25316, 
    24727, 23972,
  26844, 26811, 26692, 26754, 26503, 25481, 23889, 23090, 22508, 22434, 
    22760, 23418, 24276, 25363, 26268, 27110, 27097, 26112, 25641, 25208, 
    24572, 23917,
  26786, 26752, 26676, 26745, 26535, 25425, 23913, 23071, 22517, 22551, 
    22760, 23298, 24189, 25541, 26388, 27109, 26873, 25960, 25466, 25075, 
    24546, 23910,
  26781, 26791, 26894, 26844, 26534, 25437, 23945, 23040, 22514, 22448, 
    22742, 23360, 24139, 25339, 26363, 27169, 26837, 25903, 25504, 25099, 
    24519, 23956,
  26793, 26846, 26921, 26915, 26560, 25423, 23958, 23096, 22574, 22522, 
    22813, 23290, 24203, 25436, 26537, 27166, 26710, 25815, 25453, 25060, 
    24500, 23903,
  26777, 26834, 26797, 26863, 26491, 25458, 23932, 23102, 22580, 22502, 
    22812, 23320, 24164, 25301, 26344, 27046, 26446, 25831, 25457, 25070, 
    24468, 24012,
  26702, 26740, 26653, 26674, 26417, 25454, 24006, 23083, 22577, 22498, 
    22823, 23295, 24209, 25176, 26006, 26778, 26284, 25785, 25420, 25084, 
    24494, 23971,
  26568, 26596, 26544, 26606, 26373, 25431, 24028, 23126, 22584, 22521, 
    22882, 23342, 24253, 25348, 26499, 26570, 26291, 25847, 25503, 25113, 
    24487, 24004,
  26425, 26452, 26438, 26481, 26310, 25344, 23993, 23147, 22601, 22543, 
    22734, 23310, 24179, 25285, 26584, 26461, 26237, 25897, 25557, 25164, 
    24544, 23904,
  26316, 26355, 26395, 26454, 26257, 25405, 24030, 23191, 22643, 22533, 
    22802, 23357, 24122, 25443, 26459, 26401, 26020, 25863, 25576, 25202, 
    24588, 24079,
  26253, 26307, 26418, 26441, 26196, 25331, 24031, 23158, 22659, 22580, 
    22840, 23273, 24145, 25397, 26271, 26391, 25972, 25827, 25549, 25197, 
    24626, 24051,
  26215, 26283, 26395, 26444, 26229, 25372, 24016, 23184, 22637, 22491, 
    22736, 23257, 24048, 25306, 26313, 26328, 26026, 25891, 25557, 25171, 
    24658, 24073,
  26160, 26231, 26301, 26363, 26154, 25321, 23985, 23211, 22652, 22517, 
    22821, 23308, 24131, 25346, 26216, 26267, 26006, 25853, 25507, 25121, 
    24651, 24013,
  26029, 26112, 26225, 26338, 26138, 25321, 24030, 23197, 22666, 22556, 
    22782, 23327, 24065, 25360, 26566, 26141, 25950, 25769, 25479, 25107, 
    24600, 23954,
  26122, 26078, 26412, 26467, 26118, 25318, 24026, 23091, 22553, 22533, 
    22792, 23219, 24141, 25237, 26012, 26170, 25810, 25671, 25418, 25070, 
    24483, 23954,
  25485, 25580, 25955, 26135, 26087, 25350, 24011, 23255, 22646, 22612, 
    22813, 23429, 24314, 25523, 26635, 25854, 25700, 25822, 25548, 25238, 
    24589, 24064,
  25152, 25232, 25922, 26140, 26028, 25329, 24059, 23235, 22662, 22563, 
    22839, 23306, 24178, 25408, 26249, 25807, 25834, 25887, 25582, 25238, 
    24673, 24113,
  25180, 25119, 26207, 26326, 26057, 25265, 24019, 23132, 22629, 22547, 
    22712, 23244, 24089, 25244, 26191, 25950, 25660, 25735, 25521, 25194, 
    24560, 24075,
  25022, 24939, 26194, 26270, 26032, 25276, 24016, 23177, 22588, 22562, 
    22826, 23351, 24197, 25503, 26489, 25910, 25349, 25591, 25480, 25163, 
    24521, 23980,
  24710, 24729, 25703, 26007, 26048, 25323, 24070, 23236, 22694, 22593, 
    22851, 23354, 24180, 25270, 26300, 25663, 25659, 25785, 25520, 25203, 
    24692, 23986,
  24842, 24824, 25729, 26031, 26004, 25296, 24039, 23238, 22718, 22607, 
    22818, 23328, 24277, 25201, 26422, 25642, 25634, 25625, 25428, 25110, 
    24590, 24047,
  25034, 25008, 25778, 26059, 25990, 25284, 24005, 23228, 22706, 22592, 
    22800, 23328, 24187, 25186, 26299, 25672, 25672, 25681, 25453, 25243, 
    24712, 24017,
  25522, 25376, 26116, 26306, 26089, 25318, 23974, 23153, 22620, 22539, 
    22803, 23257, 24076, 25209, 26390, 25903, 25629, 25656, 25507, 25175, 
    24649, 24081,
  25701, 25559, 26192, 26340, 26141, 25310, 24012, 23147, 22641, 22532, 
    22803, 23295, 24284, 25258, 26070, 25984, 25679, 25634, 25445, 25175, 
    24591, 24215,
  25546, 25508, 25943, 26168, 26119, 25343, 24051, 23242, 22735, 22560, 
    22843, 23317, 24027, 25216, 26314, 25857, 25825, 25766, 25587, 25338, 
    24671, 24188,
  25563, 25497, 25974, 26231, 26150, 25353, 24089, 23232, 22715, 22632, 
    22840, 23416, 24040, 25493, 26161, 25932, 25732, 25687, 25502, 25216, 
    24690, 24161,
  25438, 25374, 25932, 26194, 26107, 25343, 24018, 23256, 22793, 22560, 
    22879, 23317, 24269, 25071, 26084, 25907, 25557, 25539, 25451, 25318, 
    24695, 24128,
  25461, 25300, 26057, 26249, 26085, 25279, 23984, 23141, 22714, 22536, 
    22843, 23249, 24091, 25146, 26170, 25872, 25442, 25469, 25355, 25082, 
    24521, 24041,
  25073, 24945, 25834, 26120, 26032, 25251, 24044, 23129, 22644, 22596, 
    22794, 23287, 24091, 25398, 26584, 25585, 25610, 25497, 25293, 25088, 
    24560, 24047,
  24628, 24505, 25641, 26044, 26001, 25245, 23984, 23144, 22679, 22567, 
    22829, 23234, 24044, 25361, 26545, 25494, 25809, 25570, 25383, 25014, 
    24585, 24014,
  23896, 23903, 25274, 25781, 25970, 25287, 24009, 23199, 22771, 22590, 
    22939, 23375, 24234, 25414, 26426, 25215, 26094, 25806, 25502, 25254, 
    24722, 24095,
  23557, 23576, 25115, 25712, 25946, 25259, 24010, 23231, 22743, 22669, 
    22899, 23416, 24190, 25337, 26407, 25162, 26487, 26237, 25686, 25268, 
    24620, 24109,
  23473, 23521, 25085, 25727, 25931, 25305, 24035, 23234, 22715, 22663, 
    22920, 23386, 24235, 25314, 26334, 25107, 26689, 26401, 25825, 25325, 
    24646, 24124,
  23771, 23873, 25131, 25743, 25943, 25273, 24009, 23250, 22760, 22652, 
    22920, 23265, 24306, 25416, 26645, 25074, 26675, 26479, 25866, 25374, 
    24710, 24204,
  24462, 24604, 25457, 25893, 26012, 25309, 24013, 23203, 22731, 22730, 
    22786, 23433, 24250, 25317, 26322, 25392, 26606, 26548, 25969, 25369, 
    24763, 24097,
  25408, 25555, 26160, 26360, 26196, 25309, 23966, 23234, 22765, 22707, 
    22806, 23423, 24222, 25159, 26379, 26324, 27169, 26741, 26056, 25430, 
    24726, 24185,
  26346, 26493, 26879, 26838, 26416, 25355, 23945, 23208, 22784, 22681, 
    22884, 23362, 24282, 25350, 26438, 27217, 27652, 26868, 26132, 25507, 
    24830, 24193,
  27048, 27219, 27040, 26940, 26407, 25385, 23987, 23268, 22790, 22742, 
    22924, 23396, 24324, 25276, 26491, 27448, 27734, 27025, 26287, 25607, 
    24882, 24224,
  27420, 27631, 27109, 26944, 26439, 25322, 23929, 23190, 22829, 22647, 
    22926, 23378, 24331, 25542, 26433, 27435, 27752, 27066, 26376, 25707, 
    24907, 24373,
  27492, 27738, 27013, 26904, 26378, 25336, 23957, 23166, 22743, 22783, 
    22960, 23426, 24312, 25536, 26484, 27391, 27746, 27095, 26411, 25693, 
    24965, 24379,
  27359, 27596, 26967, 26893, 26399, 25271, 23909, 23195, 22776, 22701, 
    22983, 23392, 24214, 25541, 26596, 27411, 27657, 27050, 26345, 25687, 
    24890, 24320,
  27081, 27253, 26934, 26827, 26324, 25322, 23949, 23202, 22768, 22784, 
    23020, 23444, 24360, 25477, 26450, 27331, 27600, 27021, 26362, 25718, 
    24916, 24299,
  26626, 26722, 26935, 26769, 26289, 25268, 23915, 23187, 22775, 22761, 
    22952, 23484, 24335, 25320, 26687, 27305, 27581, 27003, 26382, 25639, 
    24917, 24389,
  25941, 26013, 26825, 26728, 26265, 25201, 23887, 23195, 22805, 22781, 
    22957, 23446, 24176, 25596, 26557, 27274, 27659, 27041, 26437, 25742, 
    24969, 24317,
  25064, 25175, 26431, 26478, 26179, 25155, 23848, 23187, 22813, 22810, 
    22929, 23427, 24255, 25494, 26637, 27091, 27633, 26985, 26413, 25808, 
    24989, 24218,
  24120, 24315, 25734, 26047, 25962, 25081, 23821, 23174, 22855, 22815, 
    22982, 23408, 24309, 25298, 26547, 26487, 27474, 26918, 26400, 25804, 
    25120, 24360,
  23236, 23511, 24955, 25600, 25775, 25005, 23794, 23164, 22824, 22790, 
    23001, 23488, 24317, 25541, 26780, 25650, 27017, 26967, 26464, 25919, 
    25171, 24384,
  22392, 22733, 24631, 25419, 25685, 25007, 23809, 23157, 22846, 22841, 
    22996, 23423, 24379, 25616, 26344, 25253, 26872, 26913, 26442, 25895, 
    25237, 24607,
  21485, 21864, 24475, 25295, 25610, 24943, 23775, 23152, 22826, 22799, 
    22961, 23494, 24410, 25592, 26984, 24752, 26751, 26918, 26503, 26029, 
    25346, 24527,
  20515, 20904, 24067, 25071, 25531, 24882, 23782, 23162, 22868, 22832, 
    23035, 23553, 24547, 25590, 26874, 23773, 25878, 26844, 26503, 26020, 
    25349, 24655,
  19764, 20089, 23684, 24835, 25437, 24846, 23729, 23128, 22844, 22849, 
    23039, 23479, 24371, 25598, 26602, 23125, 26096, 26864, 26524, 26101, 
    25271, 24705,
  19596, 19802, 23099, 24518, 25301, 24784, 23725, 23154, 22845, 22874, 
    23069, 23517, 24460, 25662, 26850, 22407, 25288, 26768, 26462, 26048, 
    25286, 24636,
  20158, 20216, 23519, 24799, 25393, 24764, 23668, 23149, 22887, 22889, 
    23088, 23476, 24459, 25611, 26620, 23064, 25718, 26809, 26452, 25969, 
    25288, 24631,
  21121, 21088, 25176, 25721, 25687, 24854, 23629, 23081, 22868, 22890, 
    23109, 23537, 24439, 25667, 26706, 25318, 27093, 26942, 26461, 25971, 
    25316, 24592,
  21916, 21864, 25785, 26042, 25787, 24840, 23631, 23105, 22929, 22872, 
    23090, 23625, 24518, 25619, 26458, 26447, 27495, 26944, 26407, 25929, 
    25215, 24613,
  22081, 22123, 25163, 25685, 25621, 24713, 23592, 23125, 22866, 22886, 
    23006, 23524, 24397, 25593, 26620, 25816, 27186, 26856, 26341, 25881, 
    25262, 24635,
  21632, 21794, 24191, 25174, 25418, 24657, 23608, 23103, 22862, 22896, 
    22979, 23531, 24441, 25698, 27244, 24634, 26453, 26722, 26296, 25784, 
    25142, 24576,
  20920, 21182, 23562, 24809, 25258, 24597, 23547, 23090, 22904, 22893, 
    23079, 23646, 24418, 25531, 26426, 23629, 25907, 26681, 26269, 25798, 
    25129, 24664,
  20343, 20647, 23279, 24698, 25232, 24544, 23510, 23101, 22854, 22947, 
    23102, 23603, 24548, 25882, 26650, 23101, 25700, 26615, 26235, 25828, 
    25154, 24504,
  20073, 20392, 23175, 24648, 25195, 24546, 23452, 23022, 22867, 22936, 
    23084, 23631, 24522, 25910, 26991, 22758, 25669, 26561, 26194, 25754, 
    25092, 24486,
  20134, 20428, 23326, 24697, 25171, 24503, 23415, 23040, 22910, 22847, 
    23112, 23614, 24625, 25988, 26878, 22532, 25646, 26525, 26241, 25748, 
    25073, 24467,
  20467, 20715, 23721, 24916, 25230, 24475, 23397, 23016, 22926, 22905, 
    23077, 23698, 24645, 25900, 27097, 22524, 25797, 26576, 26164, 25771, 
    25015, 24461,
  21012, 21199, 24314, 25136, 25286, 24440, 23388, 23062, 22912, 22978, 
    23132, 23687, 24736, 25884, 27041, 23126, 26023, 26547, 26176, 25801, 
    25119, 24608,
  21620, 21746, 24871, 25399, 25299, 24325, 23365, 23020, 22895, 23010, 
    23232, 23788, 24539, 25969, 26750, 23790, 26214, 26536, 26212, 25776, 
    25107, 24622,
  22000, 22093, 25149, 25544, 25313, 24281, 23332, 23022, 22912, 23052, 
    23142, 23714, 24792, 25894, 27048, 24034, 26272, 26563, 26200, 25865, 
    25261, 24515,
  21848, 21937, 25263, 25585, 25295, 24257, 23328, 23039, 22906, 22964, 
    23255, 23667, 24784, 25996, 26965, 24242, 26312, 26554, 26164, 25825, 
    25181, 24557,
  21125, 21231, 25179, 25626, 25271, 24228, 23295, 22993, 22956, 22977, 
    23160, 23789, 24849, 25944, 26997, 24260, 26456, 26592, 26132, 25724, 
    24973, 24499,
  20154, 20205, 24847, 25477, 25162, 24157, 23241, 23012, 22919, 23016, 
    23243, 23716, 24744, 26037, 27118, 23475, 26554, 26520, 26164, 25658, 
    24974, 24429,
  19417, 19234, 24675, 25392, 25087, 24097, 23167, 22981, 22899, 23015, 
    23246, 23886, 25080, 26346, 26909, 22601, 26314, 26496, 25985, 25506, 
    24939, 24325,
  19040, 18543, 25008, 25453, 25056, 23995, 23119, 22950, 22912, 23046, 
    23328, 23850, 24801, 26332, 27132, 22758, 26411, 26362, 25975, 25477, 
    24795, 24221,
  18957, 18291, 25219, 25552, 25000, 23929, 23066, 22924, 22911, 23022, 
    23257, 23828, 24982, 26292, 26863, 23028, 26283, 26250, 25721, 25187, 
    24471, 23835,
  28109, 28109, 27969, 27284, 25891, 24144, 22692, 22267, 22128, 22498, 
    22969, 23600, 24646, 25750, 26964, 28618, 28959, 28075, 27453, 26769, 
    25822, 24745,
  28097, 28099, 28049, 27359, 26022, 24336, 22858, 22323, 22203, 22560, 
    22911, 23632, 24705, 25990, 26957, 28573, 29019, 27964, 27386, 26681, 
    25797, 24618,
  28063, 28085, 27994, 27397, 26121, 24400, 22889, 22326, 22176, 22526, 
    22848, 23587, 24683, 25771, 26791, 28533, 28947, 27916, 27284, 26662, 
    25741, 24725,
  27977, 28051, 27918, 27390, 26162, 24504, 22934, 22371, 22192, 22489, 
    22910, 23566, 24428, 25853, 26887, 28403, 28775, 27777, 27142, 26650, 
    25766, 24692,
  27923, 28050, 27840, 27335, 26225, 24625, 23009, 22419, 22186, 22500, 
    22858, 23510, 24419, 25837, 26975, 28232, 28681, 27738, 27094, 26544, 
    25659, 24730,
  27874, 28044, 27690, 27362, 26319, 24667, 23097, 22486, 22224, 22501, 
    22961, 23504, 24617, 25944, 26574, 28100, 28561, 27712, 27089, 26438, 
    25512, 24536,
  27841, 28014, 27696, 27351, 26324, 24753, 23154, 22466, 22233, 22457, 
    22854, 23599, 24414, 25716, 26678, 28084, 28587, 27801, 27066, 26365, 
    25417, 24436,
  27847, 27995, 27722, 27429, 26436, 24838, 23235, 22535, 22212, 22478, 
    22911, 23486, 24397, 25859, 26700, 28159, 28647, 27722, 27037, 26251, 
    25175, 24247,
  27881, 28008, 27865, 27522, 26513, 24913, 23280, 22554, 22223, 22524, 
    22879, 23565, 24393, 25672, 26350, 28250, 28760, 27782, 26979, 26153, 
    25157, 24207,
  27887, 28015, 27860, 27537, 26594, 24973, 23403, 22634, 22240, 22535, 
    22871, 23401, 24438, 25549, 26837, 28315, 28822, 27778, 26922, 26122, 
    25048, 24202,
  27831, 27967, 27826, 27535, 26591, 25085, 23391, 22648, 22264, 22494, 
    22808, 23434, 24368, 25550, 26579, 28256, 28749, 27735, 26892, 26159, 
    25028, 24100,
  27737, 27878, 27753, 27474, 26644, 25096, 23440, 22687, 22288, 22454, 
    22870, 23401, 24440, 25389, 26979, 28137, 28626, 27681, 26862, 26031, 
    25059, 24219,
  27642, 27787, 27634, 27404, 26700, 25125, 23511, 22743, 22323, 22422, 
    22833, 23418, 24397, 25629, 26451, 27957, 28470, 27438, 26700, 25878, 
    25044, 24164,
  27588, 27710, 27501, 27319, 26568, 25181, 23588, 22786, 22357, 22510, 
    22784, 23376, 24325, 25638, 26918, 27893, 28249, 27194, 26497, 25764, 
    24819, 24182,
  27562, 27657, 27413, 27270, 26606, 25183, 23543, 22782, 22327, 22421, 
    22803, 23408, 24442, 25591, 26560, 27776, 27978, 26818, 26094, 25464, 
    24745, 24058,
  27544, 27621, 27315, 27157, 26537, 25158, 23616, 22734, 22356, 22492, 
    22838, 23317, 24389, 25535, 26237, 27610, 27511, 26412, 25835, 25293, 
    24725, 24049,
  27516, 27604, 27189, 27117, 26479, 25221, 23634, 22862, 22381, 22468, 
    22826, 23384, 24281, 25517, 26344, 27277, 26887, 26140, 25704, 25230, 
    24614, 24054,
  27490, 27596, 27143, 27068, 26497, 25235, 23662, 22829, 22386, 22507, 
    22831, 23387, 24314, 25365, 26628, 27057, 25985, 25813, 25622, 25260, 
    24728, 24186,
  27461, 27581, 27208, 27094, 26581, 25265, 23720, 22890, 22389, 22466, 
    22825, 23468, 24282, 25607, 26546, 27197, 26298, 25972, 25753, 25326, 
    24694, 24218,
  27432, 27547, 27234, 27147, 26629, 25343, 23721, 22918, 22406, 22396, 
    22865, 23301, 24308, 25617, 26765, 27400, 26863, 26225, 25807, 25332, 
    24746, 24318,
  27405, 27510, 27214, 27207, 26649, 25373, 23801, 22904, 22446, 22567, 
    22772, 23375, 24227, 25350, 26295, 27434, 27401, 26412, 25865, 25328, 
    24796, 24211,
  27390, 27470, 27175, 27200, 26631, 25393, 23836, 22953, 22509, 22491, 
    22776, 23411, 24224, 25621, 26428, 27463, 27496, 26476, 25884, 25341, 
    24776, 24231,
  27355, 27408, 27220, 27179, 26590, 25403, 23846, 22964, 22499, 22488, 
    22899, 23312, 24382, 25621, 26704, 27554, 27362, 26484, 25866, 25383, 
    24726, 24042,
  27250, 27301, 27148, 27081, 26598, 25404, 23823, 22986, 22476, 22484, 
    22882, 23333, 24353, 25632, 26506, 27575, 27357, 26466, 25771, 25245, 
    24731, 24088,
  27089, 27148, 26935, 26970, 26550, 25380, 23854, 23017, 22484, 22544, 
    22801, 23352, 24379, 25271, 26427, 27376, 27295, 26340, 25743, 25146, 
    24589, 24046,
  26951, 27002, 26625, 26796, 26436, 25378, 23891, 23030, 22518, 22485, 
    22832, 23376, 24280, 25558, 26631, 27163, 27018, 26106, 25666, 25212, 
    24573, 23956,
  26895, 26923, 26716, 26873, 26488, 25412, 23930, 23056, 22515, 22525, 
    22818, 23321, 24371, 25208, 26462, 27113, 26964, 26084, 25622, 25104, 
    24534, 23961,
  26908, 26943, 26918, 26941, 26518, 25407, 23902, 23039, 22539, 22562, 
    22909, 23358, 24312, 25276, 26690, 27281, 26882, 26062, 25515, 25096, 
    24450, 23921,
  26939, 27017, 26959, 26972, 26509, 25460, 23965, 23050, 22576, 22545, 
    22834, 23344, 24078, 25485, 26497, 27318, 26841, 25969, 25497, 25063, 
    24481, 23867,
  26941, 27056, 26981, 26914, 26472, 25447, 23957, 23085, 22576, 22493, 
    22883, 23376, 24268, 25301, 26753, 27293, 26838, 25953, 25488, 25118, 
    24449, 23847,
  26885, 26989, 26853, 26854, 26444, 25411, 23983, 23124, 22584, 22473, 
    22872, 23329, 24223, 25367, 26537, 27025, 26656, 25954, 25575, 25060, 
    24544, 23916,
  26756, 26833, 26632, 26662, 26334, 25446, 24018, 23098, 22599, 22556, 
    22882, 23343, 24145, 25342, 26610, 26638, 26244, 25815, 25524, 25073, 
    24532, 24043,
  26880, 26835, 26810, 26747, 26334, 25387, 23957, 23055, 22541, 22511, 
    22868, 23326, 24196, 25371, 26185, 26585, 25690, 25528, 25371, 25048, 
    24477, 24047,
  26683, 26649, 26726, 26642, 26271, 25373, 23998, 23058, 22570, 22551, 
    22757, 23324, 24174, 25259, 26454, 26429, 25397, 25412, 25281, 25104, 
    24535, 23933,
  26530, 26513, 26751, 26564, 26257, 25322, 23967, 23122, 22541, 22525, 
    22808, 23270, 24258, 25233, 26404, 26346, 25328, 25441, 25343, 24992, 
    24426, 23973,
  26447, 26429, 26682, 26574, 26188, 25278, 23984, 23105, 22529, 22508, 
    22802, 23338, 24275, 25464, 26270, 26335, 25434, 25412, 25239, 24911, 
    24477, 23959,
  26413, 26378, 26709, 26596, 26210, 25362, 24015, 23110, 22573, 22522, 
    22817, 23316, 24124, 25084, 26444, 26313, 25639, 25571, 25350, 25010, 
    24547, 24006,
  26368, 26322, 26650, 26550, 26162, 25325, 24012, 23119, 22573, 22530, 
    22856, 23290, 24208, 25322, 26487, 26226, 25757, 25621, 25446, 25041, 
    24540, 24086,
  26241, 26207, 26524, 26509, 26147, 25314, 24005, 23125, 22623, 22487, 
    22760, 23341, 24163, 25161, 26360, 26090, 25496, 25549, 25426, 25109, 
    24598, 24066,
  25995, 25979, 26439, 26415, 26162, 25297, 23983, 23077, 22590, 22596, 
    22805, 23318, 24102, 25298, 26328, 26035, 25409, 25527, 25446, 25060, 
    24579, 24046,
  25646, 25637, 26224, 26329, 26159, 25339, 24049, 23157, 22640, 22513, 
    22785, 23338, 24252, 25240, 26560, 26007, 25770, 25671, 25467, 25072, 
    24560, 24032,
  24943, 25059, 25831, 26050, 26020, 25272, 24065, 23192, 22664, 22569, 
    22784, 23298, 24178, 25357, 26353, 25661, 25719, 25815, 25575, 25171, 
    24615, 24090,
  24906, 24881, 26082, 26194, 26064, 25291, 24015, 23172, 22616, 22550, 
    22802, 23315, 24195, 25280, 26185, 25804, 25284, 25584, 25405, 25059, 
    24496, 24045,
  24681, 24633, 25979, 26140, 26035, 25302, 24011, 23130, 22625, 22642, 
    22776, 23251, 24287, 25333, 26487, 25765, 25576, 25628, 25481, 25134, 
    24597, 23991,
  24320, 24364, 25573, 25958, 26049, 25335, 24027, 23231, 22733, 22601, 
    22840, 23340, 24249, 25329, 26066, 25499, 25675, 25699, 25472, 25217, 
    24590, 24044,
  24427, 24419, 25643, 25947, 26013, 25316, 24121, 23254, 22731, 22615, 
    22877, 23352, 24072, 25547, 26677, 25465, 25376, 25546, 25428, 25149, 
    24692, 24090,
  24905, 24740, 25957, 26143, 26053, 25291, 24029, 23166, 22710, 22598, 
    22816, 23315, 24153, 25303, 26419, 25709, 25290, 25440, 25301, 25134, 
    24648, 24139,
  25110, 24956, 26110, 26224, 26110, 25269, 24004, 23169, 22651, 22541, 
    22842, 23203, 24017, 25401, 26197, 25782, 25134, 25281, 25204, 25040, 
    24489, 24099,
  25018, 25008, 25929, 26137, 26079, 25351, 24096, 23268, 22758, 22618, 
    22867, 23368, 24160, 25230, 26390, 25740, 25457, 25493, 25376, 25118, 
    24671, 24126,
  25448, 25282, 26242, 26388, 26153, 25328, 24022, 23160, 22713, 22559, 
    22790, 23206, 24116, 25261, 26435, 26026, 25545, 25483, 25383, 25078, 
    24470, 24092,
  25486, 25278, 26191, 26321, 26104, 25347, 24018, 23145, 22684, 22544, 
    22825, 23299, 24072, 25254, 26410, 25904, 25358, 25361, 25314, 25096, 
    24546, 24052,
  25359, 25133, 26117, 26262, 26160, 25291, 24015, 23175, 22689, 22587, 
    22754, 23373, 24185, 25203, 26381, 25868, 25496, 25491, 25398, 25072, 
    24540, 24052,
  24751, 24680, 25593, 26049, 26051, 25354, 24062, 23289, 22765, 22651, 
    22899, 23358, 24212, 25264, 26575, 25552, 25985, 25836, 25592, 25240, 
    24696, 24153,
  24590, 24402, 25772, 26046, 26067, 25305, 24053, 23181, 22701, 22653, 
    22856, 23376, 24166, 25201, 26465, 25554, 26112, 25787, 25459, 25153, 
    24630, 24039,
  24065, 23888, 25613, 25971, 26018, 25249, 24067, 23175, 22681, 22565, 
    22865, 23376, 24059, 25247, 26173, 25411, 26119, 25888, 25543, 25066, 
    24508, 24153,
  23271, 23248, 25146, 25707, 25916, 25286, 24043, 23253, 22801, 22707, 
    22938, 23296, 24201, 25312, 26300, 25105, 26453, 26203, 25731, 25274, 
    24735, 24180,
  22901, 22912, 24749, 25487, 25869, 25279, 24057, 23274, 22809, 22680, 
    22827, 23383, 24252, 25491, 26465, 24799, 26515, 26325, 25812, 25307, 
    24690, 24247,
  22801, 22849, 24678, 25470, 25824, 25269, 24065, 23262, 22779, 22691, 
    22942, 23401, 24089, 25343, 26627, 24614, 26407, 26379, 25812, 25201, 
    24633, 24108,
  23084, 23177, 24844, 25543, 25857, 25294, 23984, 23222, 22755, 22692, 
    22876, 23404, 24173, 25408, 26638, 24781, 26584, 26487, 25963, 25295, 
    24672, 24135,
  23768, 23881, 25115, 25744, 25960, 25299, 24019, 23278, 22833, 22776, 
    22901, 23354, 24320, 25355, 26175, 24981, 26647, 26635, 26031, 25428, 
    24711, 24168,
  24737, 24832, 25797, 26160, 26156, 25305, 24013, 23232, 22790, 22710, 
    22958, 23395, 24134, 25552, 26335, 25788, 26874, 26857, 26181, 25550, 
    24822, 24257,
  25736, 25809, 26675, 26726, 26346, 25362, 23996, 23220, 22789, 22755, 
    22962, 23326, 24228, 25318, 26263, 26923, 27656, 26882, 26217, 25608, 
    24817, 24231,
  26514, 26600, 27095, 26898, 26434, 25335, 23970, 23201, 22809, 22716, 
    22917, 23385, 24246, 25417, 26535, 27380, 27813, 27018, 26253, 25603, 
    24869, 24275,
  26935, 27061, 27048, 26928, 26416, 25342, 23951, 23272, 22795, 22721, 
    23074, 23385, 24129, 25338, 26388, 27395, 27706, 27016, 26245, 25547, 
    24870, 24317,
  26986, 27164, 27015, 26899, 26372, 25300, 23991, 23214, 22798, 22754, 
    23011, 23377, 24205, 25449, 26114, 27332, 27656, 26995, 26336, 25683, 
    24934, 24365,
  26742, 26940, 26992, 26866, 26342, 25300, 23922, 23242, 22815, 22793, 
    22908, 23409, 24197, 25290, 26282, 27298, 27587, 27029, 26373, 25715, 
    24985, 24345,
  26278, 26440, 26906, 26826, 26306, 25267, 23954, 23217, 22857, 22793, 
    22961, 23397, 24371, 25389, 26765, 27296, 27703, 27043, 26418, 25800, 
    25063, 24357,
  25584, 25695, 26591, 26572, 26181, 25131, 23907, 23204, 22785, 22775, 
    23005, 23476, 24304, 25421, 26661, 27192, 27709, 27076, 26515, 26008, 
    25108, 24521,
  24630, 24737, 26084, 26282, 26079, 25196, 23886, 23228, 22806, 22739, 
    23047, 23506, 24332, 25322, 26638, 26874, 27731, 27041, 26479, 25937, 
    25109, 24503,
  23482, 23645, 25365, 25806, 25830, 25069, 23854, 23159, 22812, 22842, 
    23016, 23505, 24342, 25488, 26565, 26115, 27469, 27044, 26531, 25866, 
    25180, 24504,
  22326, 22576, 24148, 25117, 25550, 24995, 23840, 23189, 22837, 22823, 
    23004, 23384, 24300, 25583, 26885, 24814, 26600, 26912, 26463, 25999, 
    25203, 24626,
  21383, 21691, 23159, 24527, 25381, 24902, 23814, 23168, 22861, 22797, 
    22994, 23424, 24349, 25600, 26614, 23593, 25558, 26751, 26520, 25983, 
    25279, 24630,
  20707, 21040, 23060, 24511, 25362, 24924, 23812, 23199, 22839, 22841, 
    23021, 23410, 24505, 25610, 26744, 23379, 25507, 26785, 26491, 26096, 
    25376, 24739,
  20182, 20520, 23711, 24904, 25476, 24891, 23736, 23179, 22846, 22819, 
    22982, 23519, 24471, 25507, 26813, 23890, 26082, 26825, 26504, 26069, 
    25276, 24598,
  19679, 20021, 24550, 25321, 25637, 24987, 23812, 23207, 22865, 22898, 
    22971, 23595, 24340, 25584, 26650, 24529, 26505, 26910, 26483, 26040, 
    25342, 24720,
  19279, 19572, 24421, 25273, 25596, 24897, 23728, 23164, 22904, 22826, 
    23032, 23411, 24448, 25766, 26641, 24478, 27040, 26944, 26490, 25947, 
    25354, 24602,
  19179, 19382, 23291, 24665, 25340, 24824, 23676, 23099, 22890, 22891, 
    23062, 23494, 24353, 25679, 26644, 23049, 25871, 26718, 26407, 25963, 
    25312, 24567,
  19496, 19593, 23034, 24575, 25311, 24776, 23670, 23156, 22892, 22875, 
    22950, 23567, 24445, 25691, 26911, 22736, 25261, 26657, 26377, 25891, 
    25332, 24803,
  20022, 20080, 24164, 25152, 25490, 24785, 23694, 23131, 22858, 22934, 
    23056, 23620, 24437, 25556, 26777, 24479, 26710, 26878, 26407, 25899, 
    25335, 24690,
  20397, 20470, 24504, 25322, 25554, 24785, 23616, 23195, 22886, 22863, 
    23066, 23480, 24462, 25837, 26608, 25214, 27187, 26859, 26380, 25888, 
    25355, 24799,
  20330, 20493, 23763, 24964, 25381, 24725, 23632, 23120, 22841, 22883, 
    23073, 23508, 24398, 25685, 26841, 24214, 26281, 26712, 26315, 25853, 
    25237, 24793,
  19904, 20153, 23088, 24511, 25204, 24616, 23603, 23104, 22872, 22930, 
    23078, 23572, 24607, 25717, 26669, 23060, 25560, 26629, 26268, 25812, 
    25206, 24654,
  19441, 19745, 22672, 24367, 25162, 24595, 23556, 23076, 22927, 22907, 
    23158, 23544, 24485, 25813, 26744, 22362, 25537, 26646, 26276, 25781, 
    25187, 24602,
  19250, 19553, 22751, 24369, 25156, 24533, 23530, 23125, 22932, 22904, 
    23098, 23556, 24460, 25785, 26834, 22160, 25585, 26608, 26208, 25744, 
    25194, 24623,
  19410, 19680, 23078, 24569, 25159, 24544, 23506, 23094, 22912, 23011, 
    23165, 23529, 24572, 25733, 26957, 22201, 25704, 26583, 26222, 25818, 
    25200, 24558,
  19861, 20059, 23581, 24801, 25226, 24527, 23462, 23051, 22906, 22876, 
    23192, 23639, 24594, 25803, 26791, 22564, 25804, 26598, 26110, 25732, 
    25054, 24552,
  20498, 20619, 24167, 25066, 25273, 24456, 23441, 23055, 22845, 22994, 
    23204, 23619, 24720, 25987, 26769, 23008, 26075, 26562, 26192, 25755, 
    25061, 24573,
  21248, 21315, 24590, 25270, 25281, 24392, 23411, 23055, 22917, 23010, 
    23171, 23542, 24574, 26022, 26853, 23481, 26101, 26548, 26184, 25710, 
    25132, 24486,
  21974, 22034, 24987, 25431, 25308, 24348, 23367, 23050, 22914, 22895, 
    23120, 23721, 24623, 25823, 26791, 23833, 26149, 26594, 26254, 25766, 
    25196, 24606,
  22410, 22516, 25196, 25527, 25299, 24310, 23331, 23014, 22934, 22964, 
    23215, 23740, 24550, 26093, 27262, 24038, 26151, 26556, 26207, 25755, 
    25229, 24667,
  22286, 22455, 25270, 25612, 25241, 24266, 23347, 23022, 22882, 23061, 
    23197, 23677, 24769, 25901, 26953, 24352, 26322, 26612, 26150, 25802, 
    25136, 24695,
  21589, 21800, 25333, 25617, 25274, 24234, 23263, 23038, 22896, 22986, 
    23167, 23725, 24675, 26068, 26754, 24476, 26454, 26557, 26078, 25626, 
    25043, 24530,
  20622, 20769, 25003, 25495, 25182, 24147, 23257, 23022, 22900, 23025, 
    23304, 23842, 24848, 26110, 26759, 23649, 26478, 26571, 26192, 25728, 
    25063, 24466,
  19819, 19721, 24758, 25418, 25093, 24078, 23239, 23007, 22962, 22991, 
    23213, 23870, 24721, 26156, 26813, 22801, 26361, 26460, 26062, 25582, 
    24990, 24396,
  19327, 18919, 25100, 25537, 25062, 24009, 23201, 22992, 22929, 23026, 
    23256, 23809, 24836, 26290, 27335, 23116, 26365, 26440, 25947, 25510, 
    24884, 24272,
  19183, 18612, 25327, 25562, 25021, 23943, 23127, 22934, 22915, 22990, 
    23303, 23863, 24953, 26514, 27292, 23372, 26386, 26294, 25825, 25306, 
    24700, 24020,
  28113, 28123, 27999, 27298, 25876, 24137, 22733, 22288, 22141, 22529, 
    22810, 23567, 24746, 25866, 26782, 28684, 28981, 28053, 27435, 26742, 
    25741, 24630,
  28101, 28111, 27978, 27387, 26018, 24317, 22806, 22340, 22170, 22576, 
    23025, 23601, 24702, 26010, 26826, 28650, 29040, 28050, 27381, 26630, 
    25734, 24669,
  28069, 28096, 28010, 27456, 26092, 24418, 22901, 22328, 22203, 22553, 
    22970, 23709, 24713, 25802, 26729, 28548, 28951, 27945, 27287, 26581, 
    25660, 24582,
  27990, 28066, 27907, 27466, 26221, 24514, 22958, 22361, 22168, 22565, 
    22937, 23674, 24589, 25800, 26479, 28477, 28741, 27835, 27172, 26556, 
    25640, 24682,
  27944, 28070, 27787, 27368, 26266, 24607, 23074, 22430, 22180, 22559, 
    22986, 23674, 24468, 25757, 26819, 28303, 28597, 27732, 27172, 26542, 
    25609, 24615,
  27892, 28064, 27769, 27368, 26299, 24613, 23090, 22453, 22215, 22507, 
    22855, 23550, 24504, 25565, 26726, 28201, 28645, 27734, 27084, 26400, 
    25487, 24574,
  27838, 28019, 27709, 27362, 26354, 24787, 23140, 22495, 22223, 22507, 
    22868, 23500, 24532, 25853, 26572, 28147, 28546, 27795, 27049, 26262, 
    25260, 24374,
  27810, 27974, 27696, 27389, 26424, 24831, 23197, 22484, 22214, 22520, 
    22911, 23498, 24501, 25705, 26572, 28138, 28619, 27750, 26992, 26188, 
    25177, 24299,
  27810, 27958, 27791, 27437, 26495, 24914, 23311, 22565, 22242, 22597, 
    22865, 23534, 24428, 25538, 26544, 28330, 28725, 27825, 27106, 26194, 
    25165, 24253,
  27797, 27953, 27754, 27457, 26518, 24989, 23329, 22538, 22271, 22459, 
    22853, 23581, 24435, 25801, 26758, 28301, 28706, 27678, 26944, 26046, 
    25075, 24174,
  27743, 27906, 27732, 27428, 26590, 25067, 23394, 22647, 22304, 22490, 
    22828, 23487, 24281, 25788, 26668, 28232, 28632, 27512, 26729, 25971, 
    25017, 24045,
  27662, 27817, 27621, 27421, 26613, 25131, 23426, 22674, 22260, 22516, 
    22804, 23485, 24373, 25437, 26584, 28110, 28424, 27501, 26658, 25954, 
    25021, 24131,
  27577, 27719, 27532, 27346, 26610, 25140, 23484, 22690, 22307, 22435, 
    22790, 23472, 24383, 25619, 26550, 27991, 28292, 27250, 26522, 25697, 
    24758, 24183,
  27528, 27643, 27413, 27293, 26563, 25146, 23525, 22746, 22300, 22534, 
    22903, 23393, 24412, 25442, 26740, 27822, 28052, 26826, 26085, 25396, 
    24705, 24027,
  27506, 27605, 27408, 27225, 26537, 25198, 23554, 22699, 22332, 22482, 
    22782, 23397, 24368, 25582, 26660, 27710, 27744, 26543, 25903, 25301, 
    24664, 24109,
  27491, 27586, 27304, 27150, 26493, 25157, 23623, 22792, 22387, 22485, 
    22878, 23463, 24271, 25618, 26883, 27472, 27551, 26390, 25756, 25186, 
    24643, 24074,
  27455, 27564, 27158, 27039, 26434, 25202, 23627, 22814, 22339, 22487, 
    22877, 23374, 24385, 25437, 26802, 27192, 26926, 26153, 25673, 25216, 
    24558, 24032,
  27408, 27525, 27041, 27031, 26468, 25178, 23659, 22849, 22379, 22468, 
    22837, 23379, 24283, 25421, 26660, 26924, 26061, 25899, 25610, 25216, 
    24678, 24117,
  27350, 27473, 27178, 27079, 26559, 25267, 23730, 22864, 22406, 22520, 
    22912, 23445, 24267, 25646, 26601, 27109, 26531, 26043, 25638, 25182, 
    24644, 24028,
  27301, 27417, 27183, 27140, 26582, 25328, 23773, 22923, 22428, 22543, 
    22876, 23369, 24330, 25390, 26428, 27393, 27116, 26131, 25630, 25238, 
    24639, 24109,
  27274, 27382, 27164, 27117, 26633, 25390, 23780, 22941, 22434, 22517, 
    22864, 23390, 24217, 25519, 26661, 27432, 27310, 26268, 25790, 25264, 
    24728, 24197,
  27275, 27364, 27240, 27151, 26678, 25411, 23818, 22917, 22456, 22467, 
    22837, 23337, 24258, 25590, 26504, 27510, 27485, 26396, 25859, 25352, 
    24721, 24229,
  27258, 27327, 27314, 27169, 26629, 25418, 23873, 22975, 22462, 22555, 
    22815, 23385, 24245, 25642, 25952, 27642, 27601, 26491, 25903, 25314, 
    24695, 24168,
  27173, 27247, 27135, 27071, 26594, 25417, 23913, 23045, 22487, 22576, 
    22801, 23449, 24226, 25508, 26546, 27548, 27453, 26414, 25807, 25306, 
    24688, 24234,
  27046, 27136, 26879, 26887, 26468, 25412, 23918, 23039, 22554, 22600, 
    22765, 23410, 24364, 25373, 26645, 27271, 27216, 26275, 25649, 25157, 
    24539, 23896,
  26962, 27056, 26790, 26812, 26424, 25337, 23874, 23059, 22509, 22498, 
    22901, 23312, 24297, 25450, 26134, 27129, 26952, 26047, 25593, 25129, 
    24498, 23975,
  26970, 27051, 26922, 26910, 26501, 25399, 23898, 23063, 22576, 22567, 
    22864, 23344, 24379, 25447, 26906, 27241, 26929, 26084, 25706, 25121, 
    24535, 23799,
  27032, 27123, 27013, 26992, 26514, 25419, 23950, 23059, 22576, 22538, 
    22829, 23416, 24286, 25553, 26749, 27376, 27066, 26177, 25703, 25225, 
    24553, 24000,
  27078, 27206, 27109, 26949, 26496, 25422, 23947, 23108, 22553, 22584, 
    22897, 23389, 24140, 25444, 26464, 27403, 27154, 26229, 25727, 25217, 
    24565, 23966,
  27067, 27215, 27019, 26874, 26460, 25386, 23957, 23132, 22566, 22492, 
    22851, 23325, 24165, 25336, 26501, 27254, 27026, 26190, 25684, 25197, 
    24584, 23959,
  26982, 27104, 26846, 26736, 26402, 25404, 23993, 23102, 22589, 22569, 
    22900, 23307, 24186, 25501, 26679, 27007, 26570, 25962, 25584, 25183, 
    24609, 24048,
  26814, 26900, 26675, 26623, 26339, 25387, 24008, 23184, 22604, 22506, 
    22876, 23357, 24071, 25393, 26354, 26697, 25854, 25626, 25395, 25109, 
    24571, 24095,
  26885, 26854, 26856, 26704, 26304, 25341, 23967, 23077, 22514, 22507, 
    22780, 23359, 24145, 25375, 26159, 26651, 25230, 25087, 25145, 24891, 
    24422, 23991,
  26620, 26611, 26734, 26659, 26301, 25360, 24057, 23065, 22543, 22553, 
    22720, 23361, 24203, 25343, 26621, 26437, 25131, 25058, 25104, 24928, 
    24441, 23931,
  26400, 26409, 26635, 26582, 26212, 25299, 24012, 23080, 22549, 22607, 
    22817, 23270, 24241, 25296, 26485, 26326, 25180, 25137, 25097, 24859, 
    24389, 23998,
  26271, 26266, 26600, 26582, 26223, 25312, 24022, 23107, 22592, 22567, 
    22856, 23297, 24137, 25212, 26539, 26273, 25349, 25267, 25152, 24890, 
    24440, 23924,
  26228, 26188, 26551, 26529, 26189, 25338, 23994, 23101, 22586, 22575, 
    22796, 23226, 24198, 25247, 26493, 26203, 25330, 25310, 25193, 24921, 
    24459, 23964,
  26208, 26146, 26660, 26543, 26185, 25296, 24008, 23104, 22557, 22523, 
    22919, 23282, 23971, 25370, 26447, 26139, 25336, 25332, 25290, 24990, 
    24580, 23957,
  25800, 25883, 26320, 26287, 26166, 25362, 24050, 23244, 22676, 22551, 
    22854, 23423, 24160, 25626, 26662, 25945, 25537, 25553, 25393, 25114, 
    24627, 24004,
  25596, 25702, 26128, 26255, 26153, 25373, 24091, 23224, 22676, 22567, 
    22822, 23385, 24273, 25462, 26432, 25933, 25924, 25743, 25511, 25114, 
    24615, 24079,
  25267, 25386, 25985, 26265, 26101, 25324, 24083, 23237, 22740, 22571, 
    22934, 23426, 24209, 25322, 26091, 25843, 25897, 25843, 25523, 25145, 
    24615, 24040,
  25175, 25159, 26237, 26343, 26140, 25312, 24046, 23180, 22647, 22589, 
    22836, 23315, 24166, 25403, 25822, 25932, 25535, 25613, 25414, 25076, 
    24484, 24145,
  24773, 24753, 26104, 26204, 26103, 25298, 24035, 23165, 22656, 22560, 
    22913, 23241, 24087, 25331, 26585, 25753, 25236, 25468, 25414, 25039, 
    24491, 24057,
  24483, 24444, 25816, 26039, 25997, 25326, 24042, 23168, 22671, 22569, 
    22782, 23251, 24205, 25218, 26415, 25632, 25092, 25309, 25241, 25014, 
    24580, 24044,
  24372, 24289, 25729, 26073, 26046, 25318, 24056, 23180, 22641, 22632, 
    22952, 23413, 24195, 25284, 26404, 25577, 25036, 25338, 25324, 25101, 
    24561, 24184,
  24431, 24295, 25816, 26089, 26054, 25332, 24056, 23194, 22688, 22597, 
    22924, 23322, 24232, 25386, 26466, 25574, 25254, 25338, 25303, 25008, 
    24528, 24117,
  24596, 24428, 25831, 26073, 26063, 25320, 24035, 23209, 22720, 22574, 
    22875, 23264, 24257, 25167, 26541, 25510, 25099, 25259, 25296, 25101, 
    24624, 24198,
  24798, 24635, 25831, 26089, 26074, 25329, 24056, 23188, 22694, 22612, 
    22935, 23266, 24198, 25451, 26495, 25491, 24881, 25194, 25269, 25120, 
    24573, 24111,
  24994, 24846, 25957, 26173, 26098, 25329, 24070, 23206, 22700, 22597, 
    22901, 23357, 24141, 25191, 26497, 25716, 25329, 25446, 25358, 25039, 
    24561, 24117,
  24859, 24831, 25828, 26113, 26119, 25377, 24057, 23283, 22757, 22668, 
    22915, 23385, 24260, 25288, 26589, 25719, 25737, 25722, 25578, 25220, 
    24736, 24224,
  24894, 24833, 25809, 26148, 26115, 25351, 24130, 23309, 22757, 22670, 
    23072, 23375, 24199, 25351, 26814, 25676, 25557, 25564, 25442, 25128, 
    24640, 24197,
  24761, 24674, 25701, 26042, 26055, 25340, 24069, 23279, 22767, 22665, 
    22968, 23421, 24187, 25409, 26749, 25542, 25768, 25669, 25454, 25250, 
    24658, 24071,
  24425, 24346, 25540, 25993, 26057, 25389, 24086, 23279, 22773, 22661, 
    22947, 23370, 24311, 25393, 26606, 25430, 25925, 25713, 25408, 25221, 
    24736, 24098,
  23909, 23851, 25313, 25851, 26000, 25349, 24077, 23283, 22763, 22666, 
    22865, 23446, 24207, 25335, 26447, 25255, 26100, 25896, 25556, 25192, 
    24723, 24084,
  23304, 23273, 25098, 25729, 25900, 25327, 24085, 23278, 22798, 22696, 
    22882, 23316, 24282, 25443, 26388, 25112, 26456, 26178, 25701, 25204, 
    24653, 24226,
  22733, 22736, 24635, 25454, 25820, 25304, 24073, 23282, 22836, 22700, 
    22909, 23423, 24311, 25283, 26772, 24691, 26606, 26325, 25774, 25310, 
    24679, 24139,
  22318, 22365, 24224, 25196, 25768, 25269, 24043, 23320, 22782, 22725, 
    22926, 23408, 24272, 25586, 26438, 24082, 26231, 26491, 25890, 25262, 
    24698, 24172,
  22173, 22247, 24251, 25182, 25738, 25281, 24051, 23304, 22786, 22647, 
    22856, 23301, 24277, 25340, 26199, 23989, 26078, 26488, 25945, 25268, 
    24647, 24147,
  22374, 22461, 24533, 25355, 25813, 25264, 24036, 23265, 22783, 22687, 
    22931, 23393, 24462, 25379, 26518, 24331, 26475, 26588, 26035, 25417, 
    24744, 24147,
  22928, 23000, 24758, 25462, 25840, 25269, 23991, 23262, 22776, 22754, 
    23032, 23410, 24295, 25609, 26410, 24646, 26531, 26758, 26090, 25463, 
    24783, 24194,
  23751, 23783, 25350, 25888, 26034, 25280, 24013, 23264, 22836, 22737, 
    22961, 23382, 24383, 25304, 26522, 25326, 26789, 26813, 26210, 25567, 
    24842, 24248,
  24631, 24638, 26216, 26425, 26182, 25316, 23979, 23216, 22776, 22728, 
    22962, 23389, 24415, 25430, 26625, 26504, 27434, 26860, 26219, 25600, 
    24876, 24243,
  25334, 25362, 26796, 26707, 26312, 25335, 23948, 23256, 22797, 22801, 
    23011, 23512, 24202, 25584, 26621, 27114, 27553, 26939, 26297, 25601, 
    24832, 24227,
  25709, 25794, 26837, 26812, 26358, 25313, 23962, 23271, 22788, 22777, 
    23018, 23512, 24254, 25342, 26499, 27240, 27584, 26944, 26282, 25676, 
    24871, 24296,
  25713, 25875, 26804, 26810, 26397, 25316, 23956, 23257, 22858, 22778, 
    22979, 23532, 24345, 25492, 26616, 27251, 27615, 27031, 26400, 25731, 
    24979, 24289,
  25402, 25622, 26736, 26688, 26281, 25265, 23963, 23268, 22812, 22798, 
    23010, 23305, 24315, 25707, 26878, 27221, 27601, 27044, 26375, 25756, 
    25018, 24296,
  24852, 25081, 26471, 26461, 26137, 25232, 23934, 23243, 22894, 22828, 
    22953, 23435, 24366, 25538, 26870, 27060, 27669, 27094, 26413, 25885, 
    25064, 24329,
  24074, 24286, 25673, 25963, 25988, 25135, 23931, 23220, 22866, 22797, 
    22956, 23442, 24226, 25640, 26371, 26338, 27381, 27032, 26490, 25920, 
    25167, 24573,
  23050, 23266, 24595, 25311, 25660, 25054, 23834, 23230, 22905, 22835, 
    22913, 23452, 24209, 25567, 26874, 25245, 26562, 26897, 26502, 26047, 
    25104, 24548,
  21848, 22101, 23682, 24770, 25474, 24986, 23846, 23205, 22831, 22765, 
    22999, 23471, 24374, 25487, 26692, 24200, 25864, 26806, 26472, 25939, 
    25277, 24602,
  20661, 20960, 22699, 24256, 25231, 24873, 23818, 23176, 22833, 22796, 
    23001, 23481, 24194, 25427, 26459, 22987, 25207, 26753, 26438, 25960, 
    25223, 24617,
  19742, 20047, 22080, 23860, 25116, 24845, 23737, 23200, 22807, 22835, 
    22960, 23449, 24332, 25632, 26797, 22068, 25055, 26657, 26440, 25938, 
    25236, 24587,
  19193, 19482, 22058, 23898, 25101, 24877, 23770, 23171, 22847, 22791, 
    23057, 23455, 24362, 25563, 26595, 21929, 24792, 26684, 26410, 25989, 
    25276, 24684,
  18912, 19197, 22787, 24312, 25265, 24864, 23767, 23161, 22880, 22852, 
    23053, 23458, 24373, 25553, 26712, 22869, 25276, 26738, 26499, 25993, 
    25354, 24717,
  18709, 19020, 23845, 24931, 25456, 24884, 23732, 23189, 22887, 22810, 
    22974, 23463, 24372, 25679, 26658, 24255, 26681, 26851, 26444, 25989, 
    25356, 24665,
  18531, 18829, 23884, 24904, 25468, 24893, 23682, 23149, 22868, 22787, 
    23006, 23500, 24332, 25547, 26720, 24373, 26824, 26907, 26458, 25903, 
    25356, 24708,
  18444, 18688, 22828, 24396, 25265, 24806, 23699, 23127, 22840, 22818, 
    23045, 23450, 24404, 25598, 26554, 22908, 25617, 26782, 26444, 25949, 
    25250, 24700,
  18537, 18706, 22483, 24207, 25193, 24729, 23670, 23181, 22893, 22908, 
    23177, 23511, 24438, 25701, 26922, 22206, 25232, 26700, 26338, 25932, 
    25226, 24600,
  18716, 18869, 22992, 24442, 25304, 24749, 23665, 23146, 22948, 22889, 
    23070, 23564, 24504, 25540, 27049, 23126, 26028, 26770, 26354, 25859, 
    25260, 24709,
  18809, 18984, 23050, 24544, 25267, 24750, 23598, 23126, 22921, 22899, 
    23109, 23594, 24462, 25578, 26868, 23389, 25864, 26772, 26286, 25843, 
    25331, 24683,
  18677, 18925, 22700, 24335, 25190, 24650, 23593, 23108, 22887, 22856, 
    23059, 23612, 24432, 25668, 26890, 22629, 25436, 26634, 26324, 25807, 
    25231, 24684,
  18446, 18747, 22400, 24224, 25107, 24595, 23582, 23109, 22901, 22917, 
    23049, 23606, 24501, 25588, 26671, 22016, 25495, 26637, 26312, 25903, 
    25251, 24726,
  18371, 18691, 22481, 24279, 25120, 24613, 23551, 23093, 22917, 22928, 
    23069, 23508, 24646, 25622, 26582, 21771, 25595, 26594, 26258, 25842, 
    25176, 24573,
  18646, 18926, 22798, 24440, 25125, 24554, 23512, 23107, 22919, 22897, 
    23137, 23648, 24617, 25878, 27099, 21921, 25680, 26557, 26217, 25755, 
    25042, 24561,
  19232, 19441, 23411, 24715, 25232, 24470, 23489, 23087, 22902, 22961, 
    23150, 23551, 24587, 25866, 26721, 22385, 25824, 26533, 26128, 25618, 
    25010, 24455,
  19994, 20103, 24114, 25047, 25271, 24525, 23468, 23068, 22949, 22983, 
    23100, 23605, 24651, 25860, 26882, 23096, 26093, 26533, 26057, 25581, 
    24998, 24423,
  20803, 20832, 24515, 25273, 25344, 24471, 23459, 23072, 22924, 22958, 
    23153, 23684, 24628, 25932, 27100, 23679, 26288, 26518, 26104, 25616, 
    25004, 24491,
  21617, 21617, 24762, 25362, 25334, 24399, 23424, 23068, 22977, 22965, 
    23170, 23684, 24636, 25866, 26884, 23887, 26290, 26540, 26082, 25684, 
    25044, 24471,
  22346, 22386, 25005, 25485, 25296, 24383, 23404, 23094, 22946, 22976, 
    23105, 23698, 24720, 25900, 26913, 23820, 26089, 26558, 26153, 25753, 
    25115, 24572,
  22773, 22905, 25226, 25616, 25312, 24339, 23390, 23060, 22951, 22965, 
    23240, 23609, 24615, 26010, 27261, 23886, 26053, 26563, 26141, 25723, 
    25224, 24585,
  22661, 22882, 25329, 25679, 25305, 24301, 23305, 23045, 22931, 22977, 
    23174, 23780, 24726, 26081, 26713, 24267, 26249, 26482, 26070, 25645, 
    25042, 24546,
  22003, 22269, 25318, 25679, 25219, 24204, 23262, 23008, 22953, 23031, 
    23107, 23864, 24788, 26207, 27007, 24531, 26529, 26520, 26081, 25518, 
    25025, 24381,
  21065, 21260, 25054, 25582, 25175, 24137, 23278, 23030, 22943, 23012, 
    23221, 23867, 24954, 26324, 27135, 23857, 26462, 26527, 26098, 25646, 
    25071, 24452,
  20222, 20183, 24878, 25493, 25129, 24112, 23232, 23037, 22975, 23016, 
    23242, 23826, 25021, 26110, 27082, 22950, 26375, 26532, 26113, 25593, 
    25023, 24468,
  19635, 19312, 25078, 25498, 25061, 24042, 23204, 22976, 22937, 22979, 
    23284, 23775, 24962, 26316, 27238, 23244, 26324, 26484, 26041, 25558, 
    24962, 24351,
  19440, 18967, 25368, 25587, 25042, 23937, 23196, 22954, 22929, 23049, 
    23354, 23881, 24891, 26239, 27196, 23555, 26320, 26322, 25860, 25373, 
    24708, 24105,
  28113, 28102, 27937, 27309, 25870, 24165, 22730, 22253, 22144, 22545, 
    22978, 23617, 24640, 25832, 26560, 28690, 29049, 27964, 27250, 26567, 
    25575, 24613,
  28102, 28096, 27997, 27349, 26016, 24300, 22820, 22324, 22141, 22558, 
    22971, 23666, 24663, 25925, 26407, 28626, 29089, 27982, 27265, 26511, 
    25490, 24359,
  28075, 28097, 28009, 27422, 26138, 24398, 22892, 22344, 22206, 22555, 
    22962, 23554, 24585, 25725, 26837, 28561, 28957, 27920, 27231, 26512, 
    25468, 24365,
  28008, 28082, 27938, 27376, 26199, 24485, 22937, 22383, 22186, 22553, 
    22954, 23555, 24668, 25809, 26537, 28449, 28864, 27745, 27125, 26449, 
    25461, 24412,
  27975, 28094, 27862, 27357, 26245, 24556, 23043, 22389, 22183, 22495, 
    22979, 23615, 24553, 25920, 26593, 28303, 28657, 27663, 27000, 26337, 
    25449, 24465,
  27925, 28083, 27744, 27395, 26300, 24676, 23080, 22454, 22215, 22526, 
    22907, 23615, 24539, 25587, 26638, 28236, 28687, 27644, 26933, 26281, 
    25251, 24284,
  27855, 28021, 27685, 27381, 26378, 24734, 23151, 22472, 22220, 22447, 
    22862, 23513, 24378, 25566, 26510, 28225, 28632, 27698, 26932, 26169, 
    25106, 24064,
  27795, 27949, 27743, 27432, 26439, 24839, 23235, 22487, 22202, 22456, 
    22868, 23513, 24576, 25560, 26526, 28201, 28637, 27725, 26999, 26156, 
    25163, 24176,
  27758, 27907, 27750, 27474, 26458, 24882, 23287, 22610, 22248, 22490, 
    22876, 23407, 24414, 25799, 26500, 28204, 28705, 27737, 26906, 26106, 
    25094, 24070,
  27718, 27883, 27759, 27470, 26491, 24976, 23310, 22604, 22253, 22458, 
    22893, 23515, 24510, 25574, 26752, 28213, 28656, 27529, 26787, 25965, 
    24992, 24231,
  27652, 27827, 27592, 27414, 26568, 25012, 23378, 22642, 22272, 22495, 
    22873, 23426, 24523, 25817, 26575, 28100, 28475, 27328, 26612, 25950, 
    25029, 24189,
  27568, 27731, 27523, 27329, 26572, 25040, 23401, 22690, 22322, 22561, 
    22860, 23467, 24228, 25609, 26678, 27956, 28318, 27259, 26500, 25804, 
    24995, 24255,
  27484, 27626, 27425, 27246, 26524, 25089, 23487, 22671, 22363, 22489, 
    22807, 23479, 24285, 25532, 26619, 27838, 28179, 26987, 26254, 25634, 
    24834, 24247,
  27436, 27554, 27351, 27204, 26501, 25115, 23484, 22727, 22297, 22479, 
    22858, 23429, 24346, 25681, 26441, 27685, 27721, 26571, 25900, 25321, 
    24762, 24037,
  27417, 27534, 27171, 27101, 26424, 25060, 23562, 22753, 22347, 22504, 
    22839, 23347, 24144, 25397, 26749, 27513, 27307, 26274, 25772, 25282, 
    24599, 24127,
  27403, 27527, 27191, 27012, 26391, 25123, 23575, 22805, 22411, 22481, 
    22835, 23379, 24313, 25412, 26623, 27343, 27207, 26185, 25646, 25179, 
    24553, 24044,
  27359, 27488, 27112, 27026, 26441, 25216, 23627, 22821, 22382, 22512, 
    22866, 23371, 24306, 25481, 26743, 27106, 27013, 26187, 25722, 25190, 
    24570, 23929,
  27293, 27406, 27078, 27025, 26463, 25200, 23704, 22859, 22396, 22476, 
    22785, 23445, 24105, 25618, 26522, 27041, 26596, 26163, 25729, 25184, 
    24550, 23987,
  27214, 27308, 27109, 27113, 26503, 25283, 23717, 22879, 22421, 22490, 
    22811, 23396, 24186, 25378, 26657, 27203, 27009, 26185, 25763, 25145, 
    24555, 23918,
  27155, 27229, 27060, 27032, 26569, 25305, 23748, 22885, 22440, 22497, 
    22773, 23280, 24257, 25345, 26822, 27287, 27040, 26041, 25597, 25044, 
    24537, 23973,
  27134, 27200, 27051, 27017, 26580, 25382, 23787, 22963, 22481, 22542, 
    22835, 23337, 24151, 25504, 26643, 27281, 27078, 26027, 25564, 25071, 
    24543, 23906,
  27150, 27207, 27200, 27109, 26607, 25394, 23808, 22989, 22497, 22492, 
    22799, 23435, 24145, 25305, 26419, 27434, 27135, 26163, 25681, 25233, 
    24574, 23965,
  27152, 27204, 27164, 27066, 26564, 25378, 23801, 23014, 22468, 22512, 
    22873, 23431, 24290, 25478, 26493, 27563, 27188, 26200, 25614, 25164, 
    24535, 23978,
  27095, 27168, 27004, 26977, 26509, 25312, 23830, 23001, 22487, 22528, 
    22832, 23485, 24220, 25295, 26781, 27381, 27109, 26151, 25616, 25093, 
    24541, 23809,
  27017, 27113, 26886, 26832, 26426, 25344, 23907, 23023, 22492, 22519, 
    22832, 23308, 24310, 25370, 26647, 27204, 26972, 26076, 25600, 25032, 
    24456, 23901,
  26991, 27099, 26847, 26863, 26439, 25318, 23884, 23060, 22556, 22572, 
    22826, 23357, 24288, 25487, 26276, 27192, 26938, 26088, 25613, 25030, 
    24485, 23891,
  27042, 27147, 27022, 26895, 26437, 25342, 23930, 23044, 22574, 22540, 
    22815, 23354, 24123, 25512, 26202, 27301, 26940, 26181, 25701, 25096, 
    24535, 23971,
  27119, 27241, 27038, 26933, 26407, 25380, 23943, 23025, 22582, 22526, 
    22846, 23279, 24153, 25373, 26460, 27315, 27071, 26289, 25746, 25156, 
    24489, 23943,
  27158, 27308, 26978, 26800, 26368, 25351, 23927, 23051, 22559, 22526, 
    22763, 23364, 24115, 25446, 26596, 27216, 27028, 26319, 25797, 25241, 
    24494, 23983,
  27133, 27286, 26853, 26720, 26363, 25343, 23950, 23088, 22601, 22508, 
    22782, 23329, 24167, 25498, 26242, 27057, 26696, 26216, 25747, 25209, 
    24545, 23916,
  27030, 27144, 26784, 26679, 26291, 25282, 23955, 23109, 22578, 22557, 
    22868, 23337, 24248, 25135, 26587, 26926, 26532, 26074, 25604, 25176, 
    24596, 23925,
  26834, 26911, 26784, 26652, 26274, 25340, 23949, 23129, 22613, 22505, 
    22856, 23370, 24069, 25310, 26416, 26761, 26494, 25985, 25672, 25133, 
    24533, 24065,
  26537, 26620, 26602, 26597, 26290, 25345, 24006, 23160, 22615, 22531, 
    22832, 23358, 24242, 25386, 26412, 26697, 26152, 25881, 25562, 25119, 
    24539, 24024,
  26190, 26301, 26490, 26556, 26254, 25345, 23978, 23145, 22598, 22532, 
    22815, 23342, 24262, 25496, 26618, 26544, 25891, 25677, 25471, 25059, 
    24539, 24045,
  25878, 26004, 26293, 26432, 26182, 25370, 24008, 23159, 22643, 22568, 
    22858, 23385, 24338, 25454, 26551, 26368, 25768, 25551, 25326, 25040, 
    24499, 24004,
  25672, 25778, 26157, 26355, 26188, 25332, 24016, 23153, 22662, 22555, 
    22841, 23280, 24279, 25283, 26306, 26163, 25440, 25427, 25318, 25010, 
    24474, 23984,
  25922, 25853, 26441, 26529, 26179, 25320, 24005, 23108, 22616, 22537, 
    22853, 23376, 24196, 25439, 26154, 26217, 25198, 25170, 25077, 24883, 
    24471, 23907,
  25927, 25827, 26500, 26507, 26253, 25320, 23991, 23131, 22601, 22586, 
    22862, 23305, 24105, 25479, 26184, 26240, 25428, 25357, 25208, 24896, 
    24491, 23994,
  25591, 25620, 26299, 26354, 26224, 25375, 24085, 23207, 22673, 22605, 
    22866, 23253, 24175, 25448, 26355, 26143, 25891, 25666, 25512, 25132, 
    24588, 24122,
  25472, 25514, 26269, 26349, 26190, 25364, 24081, 23229, 22679, 22598, 
    22890, 23232, 24293, 25320, 26401, 26189, 26017, 25841, 25525, 25132, 
    24627, 24023,
  25206, 25264, 26174, 26260, 26142, 25387, 24087, 23235, 22655, 22595, 
    22854, 23381, 24051, 25366, 26425, 26030, 25866, 25754, 25462, 25101, 
    24590, 24010,
  24821, 24886, 25997, 26209, 26097, 25351, 24085, 23298, 22763, 22664, 
    22906, 23340, 24287, 25312, 26632, 25813, 25470, 25624, 25413, 25020, 
    24571, 24046,
  24715, 24651, 26001, 26165, 26084, 25300, 24018, 23157, 22645, 22606, 
    22822, 23256, 24183, 25192, 26079, 25735, 25048, 25328, 25297, 25026, 
    24611, 24081,
  24388, 24303, 25701, 26028, 26004, 25331, 24063, 23160, 22653, 22614, 
    22858, 23334, 24171, 25334, 26409, 25505, 24699, 25061, 25152, 24945, 
    24515, 24101,
  24235, 24107, 25642, 25995, 25946, 25322, 24032, 23181, 22689, 22602, 
    22841, 23388, 24062, 25421, 26266, 25480, 24904, 25198, 25214, 25013, 
    24643, 24027,
  24260, 24084, 25823, 26063, 26001, 25295, 24067, 23204, 22691, 22640, 
    22793, 23286, 24134, 25351, 26304, 25532, 25054, 25213, 25228, 24983, 
    24579, 24094,
  24399, 24200, 25764, 26041, 26026, 25300, 24067, 23175, 22683, 22568, 
    22827, 23375, 24178, 25378, 26157, 25452, 25041, 25328, 25304, 25044, 
    24604, 24155,
  24587, 24396, 25682, 26010, 26006, 25286, 24043, 23198, 22703, 22576, 
    22864, 23324, 24188, 25264, 26257, 25343, 25203, 25343, 25345, 25051, 
    24623, 24215,
  24775, 24604, 25762, 26051, 26018, 25306, 24043, 23166, 22712, 22582, 
    22804, 23373, 24218, 25381, 26465, 25502, 25701, 25595, 25462, 25181, 
    24604, 24155,
  24921, 24749, 25828, 26114, 26060, 25320, 24039, 23187, 22709, 22620, 
    22861, 23289, 24047, 25238, 26438, 25572, 25707, 25689, 25470, 25156, 
    24592, 24155,
  24970, 24773, 25875, 26106, 26047, 25337, 24029, 23151, 22686, 22631, 
    22819, 23395, 24146, 25320, 26514, 25663, 25615, 25523, 25393, 25094, 
    24573, 24208,
  24555, 24475, 25644, 26040, 26084, 25290, 24083, 23286, 22796, 22673, 
    22877, 23329, 24193, 25327, 26409, 25549, 25853, 25644, 25489, 25199, 
    24740, 24189,
  24223, 24159, 25590, 25979, 26046, 25321, 24041, 23251, 22787, 22706, 
    22833, 23261, 24198, 25225, 26506, 25474, 26085, 25768, 25533, 25201, 
    24690, 24155,
  23689, 23663, 25227, 25754, 25941, 25292, 24040, 23264, 22830, 22694, 
    22931, 23319, 24165, 25418, 26099, 25236, 26293, 26009, 25619, 25223, 
    24646, 24196,
  23046, 23066, 24752, 25475, 25812, 25293, 24068, 23270, 22812, 22684, 
    22865, 23460, 24218, 25456, 26704, 24751, 26518, 26253, 25764, 25278, 
    24773, 24143,
  22428, 22495, 24193, 25185, 25703, 25236, 24070, 23300, 22783, 22740, 
    22960, 23344, 24309, 25436, 26606, 24090, 26343, 26394, 25857, 25291, 
    24716, 24156,
  21954, 22056, 24135, 25118, 25682, 25233, 24040, 23265, 22814, 22686, 
    22927, 23337, 24290, 25346, 26529, 23812, 26175, 26451, 25876, 25312, 
    24640, 24156,
  21698, 21798, 24084, 25096, 25647, 25225, 24066, 23268, 22862, 22747, 
    22853, 23308, 24186, 25645, 26579, 23871, 26432, 26585, 26007, 25437, 
    24780, 24191,
  21688, 21764, 24169, 25145, 25685, 25185, 23994, 23284, 22836, 22761, 
    22939, 23304, 24191, 25481, 26762, 23978, 26274, 26664, 26125, 25460, 
    24812, 24191,
  21924, 21960, 24362, 25244, 25772, 25229, 24016, 23296, 22823, 22711, 
    22966, 23399, 24251, 25524, 26630, 24195, 26412, 26668, 26146, 25432, 
    24757, 24157,
  22378, 22371, 24653, 25468, 25844, 25241, 23996, 23268, 22809, 22676, 
    22998, 23440, 24275, 25389, 26591, 24670, 26451, 26760, 26135, 25461, 
    24810, 24245,
  22922, 22906, 25282, 25826, 25951, 25242, 23979, 23253, 22899, 22779, 
    22965, 23429, 24194, 25459, 26615, 25573, 26966, 26822, 26192, 25556, 
    24856, 24179,
  23389, 23412, 25846, 26193, 26112, 25257, 23980, 23242, 22832, 22768, 
    22959, 23367, 24415, 25560, 26475, 26406, 27478, 26957, 26346, 25619, 
    24965, 24291,
  23643, 23736, 26108, 26294, 26115, 25264, 23928, 23248, 22820, 22716, 
    22926, 23407, 24371, 25329, 26339, 26663, 27545, 27006, 26435, 25707, 
    24973, 24393,
  23628, 23812, 26015, 26266, 26112, 25208, 23971, 23249, 22797, 22757, 
    23019, 23443, 24225, 25433, 26186, 26685, 27589, 27093, 26421, 25804, 
    25024, 24393,
  23377, 23644, 25637, 26060, 26007, 25180, 23890, 23254, 22839, 22771, 
    22990, 23426, 24146, 25641, 26691, 26446, 27600, 27112, 26466, 25854, 
    25112, 24493,
  22950, 23262, 25083, 25696, 25816, 25153, 23914, 23256, 22859, 22776, 
    23058, 23440, 24386, 25302, 26423, 25859, 27331, 26982, 26484, 25890, 
    25178, 24420,
  22349, 22669, 24232, 25153, 25536, 25022, 23886, 23225, 22846, 22822, 
    22927, 23412, 24284, 25679, 26679, 24666, 26421, 26827, 26435, 25925, 
    25185, 24477,
  21540, 21859, 23512, 24643, 25370, 24964, 23882, 23208, 22864, 22814, 
    22996, 23325, 24360, 25647, 26388, 23526, 25446, 26706, 26454, 25935, 
    25199, 24444,
  20552, 20873, 23078, 24385, 25252, 24910, 23829, 23253, 22916, 22817, 
    23030, 23484, 24187, 25596, 26531, 22871, 25377, 26716, 26514, 26025, 
    25264, 24600,
  19530, 19850, 22495, 24070, 25161, 24859, 23815, 23199, 22888, 22810, 
    23030, 23543, 24369, 25501, 26651, 22259, 25168, 26669, 26500, 26001, 
    25401, 24621,
  18703, 18991, 22031, 23826, 25094, 24852, 23831, 23213, 22898, 22868, 
    22931, 23502, 24283, 25607, 26555, 21698, 24830, 26654, 26454, 25962, 
    25305, 24585,
  18196, 18451, 21872, 23701, 25064, 24838, 23762, 23187, 22908, 22853, 
    23032, 23432, 24377, 25632, 26695, 21531, 24822, 26666, 26521, 25976, 
    25326, 24661,
  17960, 18212, 22030, 23871, 25103, 24774, 23743, 23194, 22863, 22911, 
    22996, 23543, 24451, 25515, 26806, 21969, 24994, 26685, 26500, 25999, 
    25392, 24741,
  17824, 18123, 22486, 24186, 25179, 24780, 23732, 23190, 22840, 22812, 
    23011, 23503, 24306, 25603, 26622, 22812, 25521, 26719, 26445, 26001, 
    25324, 24683,
  17695, 18009, 22533, 24186, 25182, 24775, 23708, 23200, 22903, 22826, 
    22947, 23474, 24404, 25613, 26893, 22824, 25651, 26702, 26438, 25928, 
    25362, 24604,
  17564, 17849, 22105, 23950, 25060, 24684, 23659, 23132, 22889, 22825, 
    23006, 23521, 24358, 25653, 26663, 22020, 25255, 26693, 26293, 25886, 
    25313, 24750,
  17498, 17720, 21970, 23919, 25059, 24720, 23657, 23147, 22840, 22873, 
    23055, 23495, 24423, 25410, 26492, 21607, 25212, 26669, 26332, 25901, 
    25371, 24778,
  17474, 17676, 22068, 23963, 25086, 24698, 23650, 23150, 22916, 22914, 
    23108, 23477, 24416, 25890, 26821, 21915, 25355, 26658, 26389, 25947, 
    25246, 24806,
  17452, 17660, 22231, 24060, 25084, 24654, 23606, 23112, 22909, 22918, 
    23117, 23581, 24432, 25819, 26968, 21977, 25340, 26632, 26321, 25810, 
    25190, 24620,
  17399, 17662, 22240, 24042, 25089, 24616, 23568, 23150, 22869, 22878, 
    23121, 23586, 24379, 25691, 26686, 21739, 25404, 26631, 26249, 25781, 
    25211, 24655,
  17460, 17761, 22304, 24125, 25092, 24566, 23554, 23160, 22921, 22914, 
    23114, 23626, 24430, 25687, 26834, 21621, 25518, 26654, 26375, 25784, 
    25200, 24636,
  17816, 18118, 22538, 24276, 25132, 24553, 23535, 23123, 22911, 22908, 
    23123, 23604, 24483, 25975, 26997, 21720, 25638, 26641, 26294, 25767, 
    25143, 24644,
  18534, 18776, 23121, 24545, 25186, 24514, 23509, 23134, 22974, 23020, 
    23155, 23673, 24571, 25692, 27119, 22099, 25642, 26554, 26176, 25704, 
    25022, 24458,
  19462, 19620, 23919, 24898, 25281, 24558, 23521, 23092, 22970, 22988, 
    23056, 23638, 24512, 25939, 26710, 22926, 25990, 26457, 26135, 25660, 
    24914, 24325,
  20406, 20469, 24485, 25211, 25323, 24477, 23456, 23081, 22975, 22962, 
    23214, 23641, 24562, 25915, 26874, 23737, 26303, 26457, 26121, 25512, 
    24806, 24320,
  21249, 21254, 24759, 25349, 25313, 24440, 23466, 23067, 22965, 23009, 
    23255, 23621, 24619, 25850, 27194, 24105, 26399, 26501, 26057, 25603, 
    24990, 24414,
  22004, 22012, 24830, 25418, 25323, 24385, 23411, 23082, 22934, 22968, 
    23142, 23665, 24523, 25944, 26950, 23951, 26320, 26588, 26110, 25671, 
    25114, 24521,
  22658, 22722, 24961, 25453, 25265, 24357, 23360, 23024, 22940, 23014, 
    23245, 23711, 24671, 25754, 27012, 23734, 26119, 26526, 26154, 25713, 
    25146, 24615,
  23048, 23197, 25176, 25549, 25279, 24299, 23366, 23056, 22960, 22984, 
    23198, 23670, 24699, 26138, 26725, 23803, 25959, 26596, 26210, 25709, 
    25198, 24656,
  22959, 23177, 25363, 25634, 25235, 24239, 23334, 23023, 22907, 23019, 
    23186, 23742, 24777, 26127, 26904, 24337, 26303, 26572, 26112, 25707, 
    25029, 24396,
  22369, 22614, 25459, 25710, 25245, 24223, 23287, 23027, 22959, 23082, 
    23261, 23785, 24887, 26012, 26824, 24635, 26573, 26553, 26081, 25568, 
    24967, 24425,
  21486, 21662, 25154, 25560, 25188, 24203, 23268, 23049, 22949, 23043, 
    23274, 23804, 24848, 26228, 27015, 24075, 26566, 26510, 26126, 25620, 
    24987, 24489,
  20627, 20594, 24872, 25475, 25138, 24107, 23246, 23032, 22951, 23041, 
    23310, 23899, 24990, 26234, 27340, 23121, 26404, 26501, 26100, 25493, 
    25003, 24492,
  19966, 19685, 25024, 25462, 25036, 24029, 23177, 23025, 22970, 23030, 
    23250, 23833, 24928, 26123, 26876, 23233, 26472, 26459, 26075, 25576, 
    25050, 24462,
  19727, 19314, 25279, 25504, 24986, 23942, 23162, 22996, 22956, 23028, 
    23300, 23936, 25062, 26322, 27290, 23549, 26412, 26435, 25910, 25428, 
    24841, 24329,
  28098, 28060, 28019, 27240, 25895, 24159, 22749, 22274, 22155, 22545, 
    22919, 23648, 24770, 25969, 26332, 28729, 29079, 27994, 27319, 26543, 
    25669, 24593,
  28089, 28067, 27967, 27329, 26031, 24264, 22822, 22270, 22146, 22535, 
    22832, 23573, 24429, 25816, 26782, 28613, 29057, 28028, 27403, 26605, 
    25612, 24539,
  28071, 28095, 28011, 27394, 26119, 24412, 22891, 22353, 22231, 22537, 
    22974, 23630, 24545, 25883, 26610, 28576, 29079, 28038, 27287, 26581, 
    25582, 24579,
  28018, 28103, 28000, 27397, 26186, 24490, 22950, 22430, 22209, 22518, 
    22908, 23627, 24618, 25841, 26854, 28517, 28919, 27920, 27283, 26481, 
    25600, 24579,
  27995, 28119, 27862, 27379, 26266, 24567, 23055, 22430, 22205, 22575, 
    22953, 23527, 24496, 25764, 26896, 28357, 28726, 27679, 27000, 26294, 
    25346, 24357,
  27950, 28096, 27891, 27424, 26300, 24640, 23127, 22442, 22231, 22543, 
    22951, 23560, 24635, 25721, 26682, 28295, 28699, 27661, 26904, 26232, 
    25276, 24203,
  27873, 28010, 27766, 27394, 26419, 24757, 23195, 22516, 22263, 22543, 
    22821, 23508, 24542, 25761, 26703, 28192, 28700, 27721, 27000, 26262, 
    25213, 24204,
  27790, 27907, 27721, 27450, 26460, 24822, 23234, 22567, 22254, 22490, 
    22870, 23589, 24467, 25870, 26626, 28242, 28667, 27762, 27033, 26163, 
    25188, 24289,
  27718, 27829, 27719, 27400, 26477, 24922, 23303, 22583, 22287, 22501, 
    22889, 23585, 24584, 25764, 26619, 28169, 28630, 27724, 26934, 26187, 
    25144, 24229,
  27642, 27774, 27647, 27394, 26479, 24985, 23374, 22671, 22285, 22579, 
    22987, 23599, 24453, 25704, 26850, 28107, 28488, 27547, 26800, 26101, 
    25054, 24183,
  27550, 27698, 27554, 27327, 26493, 25008, 23418, 22668, 22277, 22509, 
    22783, 23510, 24384, 25587, 26822, 27960, 28257, 27257, 26578, 25921, 
    25136, 24417,
  27456, 27593, 27435, 27237, 26532, 25037, 23460, 22681, 22289, 22549, 
    22833, 23454, 24321, 25623, 26534, 27809, 28018, 27030, 26244, 25651, 
    24975, 24268,
  27378, 27491, 27349, 27128, 26486, 25118, 23496, 22712, 22315, 22446, 
    22820, 23492, 24237, 25551, 26865, 27682, 27836, 26685, 26019, 25442, 
    24794, 24126,
  27343, 27433, 27216, 27047, 26415, 25078, 23513, 22724, 22311, 22526, 
    22859, 23351, 24387, 25610, 26640, 27482, 27446, 26370, 25844, 25260, 
    24659, 24077,
  27333, 27433, 27069, 26944, 26387, 25087, 23554, 22752, 22340, 22512, 
    22867, 23344, 24362, 25660, 26538, 27215, 27057, 26160, 25676, 25257, 
    24649, 23912,
  27317, 27432, 27010, 26928, 26358, 25115, 23587, 22810, 22416, 22498, 
    22839, 23370, 24288, 25585, 26813, 26959, 26614, 25971, 25563, 25124, 
    24527, 23943,
  27259, 27374, 27028, 26930, 26368, 25137, 23650, 22853, 22446, 22507, 
    22881, 23439, 24308, 25429, 26517, 26953, 26669, 26044, 25660, 25141, 
    24651, 24121,
  27169, 27255, 27068, 27016, 26497, 25236, 23654, 22876, 22461, 22507, 
    22909, 23394, 24302, 25471, 26984, 27131, 27062, 26331, 25818, 25315, 
    24662, 23979,
  27070, 27125, 26984, 27029, 26493, 25292, 23719, 22894, 22437, 22501, 
    22889, 23359, 24238, 25464, 26518, 27249, 27388, 26446, 25853, 25326, 
    24662, 23971,
  27007, 27033, 26761, 26797, 26435, 25293, 23709, 22887, 22430, 22554, 
    22923, 23361, 24192, 25490, 26588, 27134, 27325, 26382, 25804, 25089, 
    24585, 24039,
  26997, 27009, 26859, 26854, 26464, 25326, 23779, 22962, 22450, 22539, 
    22839, 23355, 24328, 25453, 26480, 27162, 27233, 26231, 25647, 25078, 
    24503, 23938,
  27028, 27035, 27119, 26987, 26560, 25330, 23831, 23009, 22499, 22537, 
    22868, 23376, 24199, 25571, 26328, 27418, 27122, 26099, 25619, 25041, 
    24528, 23985,
  27367, 27267, 27347, 27089, 26490, 25319, 23801, 22900, 22424, 22459, 
    22780, 23303, 24282, 25513, 26582, 27682, 26860, 25788, 25335, 24868, 
    24352, 23890,
  27030, 27071, 26910, 26879, 26485, 25372, 23864, 23048, 22512, 22519, 
    22829, 23398, 24265, 25493, 26594, 27340, 26947, 26009, 25506, 25020, 
    24424, 24009,
  27006, 27070, 26878, 26826, 26476, 25383, 23920, 23018, 22562, 22498, 
    22845, 23309, 24216, 25517, 26401, 27257, 27058, 26179, 25697, 25193, 
    24587, 23846,
  27028, 27105, 26976, 26913, 26431, 25347, 23918, 23080, 22543, 22506, 
    22810, 23414, 24142, 25492, 26641, 27304, 27168, 26343, 25828, 25211, 
    24637, 23911,
  27096, 27184, 26977, 26941, 26479, 25377, 23939, 23076, 22573, 22503, 
    22948, 23369, 24086, 25566, 26535, 27341, 27151, 26385, 25866, 25239, 
    24534, 23990,
  27157, 27277, 26982, 26819, 26336, 25335, 23924, 23075, 22607, 22551, 
    22853, 23441, 24290, 25471, 26644, 27249, 26982, 26299, 25828, 25243, 
    24590, 23936,
  27171, 27321, 26890, 26746, 26341, 25290, 23915, 23100, 22625, 22522, 
    22892, 23438, 24078, 25437, 26335, 27105, 26934, 26307, 25804, 25298, 
    24614, 24103,
  27127, 27272, 26851, 26768, 26344, 25321, 23931, 23138, 22609, 22519, 
    22849, 23284, 24314, 25398, 26739, 26988, 26788, 26268, 25801, 25272, 
    24633, 23989,
  27013, 27114, 26809, 26719, 26321, 25314, 23964, 23144, 22632, 22548, 
    22887, 23326, 24238, 25412, 26553, 26932, 26774, 26256, 25813, 25202, 
    24620, 23997,
  26795, 26864, 26712, 26686, 26281, 25325, 23979, 23178, 22574, 22479, 
    22832, 23393, 24163, 25409, 26143, 26971, 26779, 26275, 25797, 25289, 
    24678, 23997,
  26450, 26530, 26663, 26625, 26325, 25340, 23963, 23180, 22611, 22579, 
    22876, 23450, 24140, 25368, 26722, 26874, 26806, 26344, 25845, 25307, 
    24723, 24064,
  26024, 26131, 26529, 26571, 26270, 25323, 24025, 23153, 22618, 22466, 
    22779, 23456, 24212, 25478, 26728, 26790, 26738, 26242, 25816, 25258, 
    24633, 24091,
  25617, 25732, 26333, 26436, 26213, 25353, 24024, 23171, 22666, 22597, 
    22862, 23281, 24167, 25383, 26439, 26638, 26440, 26022, 25685, 25246, 
    24676, 24151,
  25323, 25417, 26051, 26262, 26175, 25365, 24046, 23197, 22697, 22598, 
    22791, 23376, 24251, 25387, 26706, 26378, 26179, 25826, 25546, 25110, 
    24594, 24037,
  25192, 25255, 25924, 26248, 26159, 25365, 24042, 23214, 22693, 22578, 
    22897, 23257, 24273, 25065, 26169, 26218, 26029, 25681, 25443, 25035, 
    24625, 24012,
  25206, 25224, 26072, 26259, 26159, 25351, 24024, 23235, 22707, 22557, 
    22837, 23318, 24252, 25325, 26462, 26179, 25897, 25679, 25407, 24935, 
    24529, 24120,
  25265, 25249, 26106, 26401, 26176, 25406, 24101, 23263, 22704, 22542, 
    22890, 23332, 24195, 25372, 26131, 26300, 26146, 25797, 25443, 25059, 
    24599, 24094,
  25250, 25220, 26198, 26319, 26189, 25362, 24038, 23240, 22669, 22572, 
    22737, 23347, 24179, 25381, 26469, 26346, 26382, 25800, 25476, 25058, 
    24594, 23969,
  25079, 25061, 26032, 26275, 26120, 25354, 24051, 23220, 22736, 22581, 
    22832, 23262, 24186, 25292, 26734, 26211, 26269, 25806, 25435, 24977, 
    24525, 24023,
  24759, 24757, 25878, 26147, 26061, 25343, 24043, 23263, 22692, 22560, 
    22865, 23318, 24176, 25412, 26613, 25961, 25979, 25769, 25461, 25058, 
    24538, 24025,
  24371, 24378, 25713, 26047, 26037, 25258, 24076, 23243, 22769, 22620, 
    22865, 23347, 24297, 25349, 26357, 25678, 25645, 25593, 25412, 25085, 
    24577, 24073,
  24356, 24207, 25703, 26016, 25985, 25253, 24024, 23189, 22664, 22521, 
    22811, 23342, 24013, 25346, 26207, 25550, 25059, 25308, 25255, 24909, 
    24489, 24081,
  24188, 23999, 25515, 25929, 25957, 25295, 24038, 23207, 22714, 22567, 
    22771, 23162, 24173, 25328, 26401, 25391, 25077, 25250, 25200, 24996, 
    24565, 24141,
  24187, 23969, 25696, 25997, 26031, 25303, 24020, 23178, 22679, 22576, 
    22845, 23378, 24227, 25176, 26241, 25438, 25152, 25308, 25255, 25026, 
    24520, 24087,
  24302, 24080, 25769, 26046, 26016, 25317, 24031, 23192, 22725, 22613, 
    22865, 23355, 24264, 25160, 26560, 25502, 25239, 25395, 25339, 25014, 
    24501, 23973,
  24471, 24267, 25650, 26010, 26013, 25252, 24031, 23210, 22661, 22584, 
    22769, 23320, 24126, 25283, 26478, 25438, 25569, 25539, 25387, 24996, 
    24609, 24100,
  24649, 24464, 25647, 25981, 26004, 25236, 24044, 23189, 22699, 22639, 
    22886, 23286, 24126, 25388, 26267, 25491, 25676, 25539, 25408, 24983, 
    24539, 24047,
  24793, 24611, 25678, 26035, 26019, 25270, 24038, 23201, 22714, 22656, 
    22774, 23357, 24092, 25260, 26117, 25455, 25588, 25510, 25408, 25045, 
    24616, 24148,
  24850, 24657, 25751, 26046, 25999, 25298, 23992, 23198, 22679, 22596, 
    22851, 23271, 24128, 25325, 26362, 25519, 25731, 25597, 25435, 25045, 
    24565, 24208,
  24460, 24403, 25534, 25923, 25979, 25276, 24044, 23283, 22778, 22661, 
    22927, 23380, 24198, 25371, 26793, 25445, 25990, 25725, 25462, 25051, 
    24624, 24195,
  24170, 24147, 25463, 25917, 26019, 25327, 24036, 23266, 22801, 22654, 
    22848, 23393, 24175, 25462, 26197, 25445, 26265, 25914, 25575, 25134, 
    24657, 24141,
  23978, 23870, 25325, 25844, 25945, 25259, 23992, 23210, 22714, 22634, 
    22894, 23254, 24272, 25164, 26476, 25188, 26285, 25973, 25587, 25077, 
    24622, 24154,
  23074, 23162, 24359, 25273, 25719, 25248, 24011, 23237, 22829, 22661, 
    22975, 23380, 24270, 25587, 26401, 24170, 26024, 26234, 25702, 25204, 
    24645, 24035,
  22451, 22585, 24142, 25074, 25651, 25225, 24003, 23268, 22832, 22656, 
    22910, 23261, 24311, 25322, 26338, 23684, 25906, 26266, 25809, 25304, 
    24658, 24148,
  21897, 22052, 24246, 25176, 25700, 25230, 24021, 23303, 22787, 22680, 
    22896, 23306, 24097, 25313, 26451, 23926, 26316, 26482, 25966, 25381, 
    24708, 24175,
  21443, 21570, 24051, 25036, 25624, 25180, 23995, 23262, 22835, 22721, 
    22923, 23314, 24265, 25393, 26626, 23829, 26201, 26595, 26029, 25362, 
    24696, 24163,
  21082, 21164, 23835, 24940, 25618, 25137, 24006, 23266, 22820, 22746, 
    22851, 23364, 24171, 25444, 26555, 23593, 25929, 26608, 26063, 25443, 
    24748, 24204,
  20830, 20869, 23965, 25041, 25641, 25176, 24011, 23275, 22831, 22728, 
    22997, 23368, 24303, 25427, 26312, 23947, 26491, 26721, 26110, 25507, 
    24749, 24271,
  20743, 20752, 23890, 24964, 25584, 25168, 23956, 23273, 22820, 22704, 
    22919, 23303, 24235, 25371, 26741, 24043, 26350, 26791, 26191, 25617, 
    24860, 24231,
  20811, 20824, 23796, 24894, 25640, 25135, 23988, 23276, 22869, 22758, 
    22935, 23393, 24285, 25308, 26222, 24112, 26353, 26817, 26316, 25663, 
    25001, 24380,
  20956, 21010, 23886, 24959, 25593, 25181, 23965, 23276, 22878, 22668, 
    22943, 23342, 24389, 25429, 26888, 24415, 26372, 26829, 26338, 25751, 
    24977, 24357,
  21084, 21194, 23881, 24953, 25581, 25119, 23961, 23236, 22849, 22747, 
    22982, 23357, 24210, 25351, 26488, 24552, 26603, 26906, 26393, 25745, 
    24965, 24332,
  21127, 21315, 23730, 24820, 25515, 25080, 23920, 23290, 22890, 22748, 
    22971, 23410, 24192, 25391, 26410, 24354, 26235, 26906, 26490, 25825, 
    25054, 24426,
  21086, 21360, 23517, 24670, 25444, 25051, 23931, 23251, 22876, 22765, 
    22952, 23388, 24343, 25550, 26581, 24009, 25879, 26847, 26438, 25850, 
    25048, 24440,
  20987, 21318, 23355, 24539, 25349, 25007, 23895, 23214, 22849, 22810, 
    23045, 23367, 24307, 25573, 26562, 23681, 25398, 26797, 26510, 25972, 
    25146, 24467,
  20789, 21140, 23259, 24471, 25279, 24978, 23836, 23221, 22874, 22773, 
    22997, 23356, 24412, 25530, 26426, 23232, 25336, 26771, 26449, 25994, 
    25196, 24516,
  20412, 20761, 23145, 24449, 25297, 24942, 23840, 23231, 22852, 22847, 
    23043, 23410, 24329, 25659, 26865, 22931, 25327, 26672, 26454, 25979, 
    25364, 24551,
  19822, 20161, 23141, 24401, 25265, 24908, 23835, 23241, 22904, 22782, 
    22849, 23469, 24206, 25591, 26585, 22918, 25400, 26697, 26445, 25995, 
    25301, 24620,
  19092, 19419, 22849, 24250, 25214, 24884, 23810, 23248, 22867, 22798, 
    22991, 23450, 24441, 25258, 26893, 22604, 25310, 26657, 26472, 25879, 
    25266, 24708,
  18399, 18693, 22482, 24059, 25135, 24880, 23764, 23206, 22842, 22851, 
    22983, 23459, 24308, 25370, 26707, 22116, 25271, 26706, 26488, 25988, 
    25317, 24699,
  17874, 18134, 22074, 23859, 25115, 24818, 23734, 23196, 22843, 22787, 
    22905, 23452, 24320, 25753, 26263, 21720, 25038, 26675, 26431, 25970, 
    25351, 24674,
  17536, 17787, 21787, 23736, 25042, 24777, 23762, 23203, 22873, 22860, 
    22992, 23460, 24398, 25371, 26501, 21532, 24918, 26665, 26458, 25950, 
    25327, 24808,
  17289, 17579, 21714, 23720, 24997, 24766, 23737, 23211, 22879, 22843, 
    23049, 23519, 24375, 25401, 26454, 21567, 24879, 26641, 26348, 25871, 
    25399, 24709,
  17064, 17376, 21737, 23801, 25015, 24744, 23699, 23146, 22867, 22873, 
    23002, 23529, 24444, 25474, 26930, 21568, 24904, 26653, 26424, 26009, 
    25381, 24765,
  16835, 17137, 21687, 23710, 25026, 24721, 23685, 23222, 22930, 22860, 
    22975, 23526, 24410, 25492, 26463, 21359, 24979, 26738, 26355, 25912, 
    25312, 24723,
  16655, 16904, 21793, 23775, 25032, 24707, 23683, 23159, 22940, 22846, 
    23051, 23511, 24477, 25499, 26743, 21284, 25154, 26656, 26338, 25801, 
    25307, 24765,
  16539, 16755, 21886, 23839, 25018, 24673, 23654, 23179, 22900, 22856, 
    23051, 23571, 24403, 25601, 26810, 21379, 25304, 26603, 26278, 25803, 
    25277, 24706,
  16516, 16712, 21942, 23979, 25051, 24662, 23639, 23162, 22937, 22863, 
    23088, 23630, 24471, 25831, 26590, 21436, 25282, 26554, 26225, 25799, 
    25201, 24754,
  16616, 16850, 22083, 24031, 25064, 24605, 23586, 23165, 22924, 22901, 
    23191, 23594, 24418, 25757, 26922, 21518, 25427, 26640, 26242, 25819, 
    25350, 24742,
  16983, 17247, 22294, 24170, 25050, 24605, 23609, 23157, 22926, 22899, 
    23115, 23535, 24516, 25725, 26787, 21593, 25535, 26635, 26188, 25810, 
    25287, 24877,
  17726, 17983, 22621, 24337, 25134, 24593, 23565, 23070, 22954, 22884, 
    23105, 23582, 24530, 25740, 27292, 21854, 25481, 26543, 26135, 25699, 
    25059, 24530,
  18798, 18983, 23445, 24703, 25265, 24559, 23549, 23122, 22982, 22927, 
    23116, 23582, 24497, 25692, 26779, 22489, 25684, 26520, 26156, 25691, 
    25028, 24490,
  19948, 20051, 24279, 25081, 25282, 24531, 23501, 23120, 22949, 22976, 
    23080, 23577, 24639, 25929, 26697, 23453, 26051, 26502, 26101, 25544, 
    24990, 24432,
  20946, 20982, 24693, 25312, 25339, 24457, 23512, 23121, 22968, 22844, 
    23116, 23621, 24518, 25759, 26804, 24071, 26226, 26517, 26079, 25544, 
    24958, 24427,
  21709, 21730, 24732, 25353, 25346, 24431, 23464, 23097, 22975, 22980, 
    23197, 23636, 24580, 26021, 26816, 24116, 26260, 26431, 26077, 25586, 
    24997, 24507,
  22328, 22380, 24690, 25361, 25302, 24441, 23444, 23099, 22942, 22929, 
    23120, 23615, 24471, 26037, 26985, 23829, 26213, 26489, 26118, 25616, 
    25068, 24601,
  22871, 22970, 24918, 25498, 25304, 24394, 23442, 23077, 22957, 22962, 
    23235, 23695, 24629, 25792, 26606, 23798, 26068, 26499, 26162, 25641, 
    25081, 24675,
  23224, 23369, 25346, 25666, 25326, 24326, 23375, 23064, 22912, 22921, 
    23202, 23665, 24679, 26150, 26789, 24187, 26144, 26575, 26210, 25723, 
    25146, 24595,
  23180, 23354, 25528, 25694, 25264, 24236, 23304, 23028, 22953, 22987, 
    23210, 23752, 24831, 26010, 26950, 24644, 26340, 26574, 26167, 25651, 
    25104, 24510,
  22685, 22871, 25550, 25703, 25229, 24201, 23286, 23026, 22997, 23021, 
    23171, 23691, 24594, 26238, 26904, 24890, 26490, 26519, 26053, 25537, 
    24921, 24291,
  21881, 22010, 25319, 25557, 25166, 24111, 23290, 22992, 22960, 23014, 
    23215, 23736, 24772, 26179, 27121, 24354, 26528, 26454, 26092, 25497, 
    24954, 24468,
  21031, 20978, 24965, 25447, 25071, 24090, 23266, 23040, 22928, 22986, 
    23345, 23857, 24721, 26260, 26891, 23274, 26435, 26416, 25969, 25512, 
    24983, 24445,
  20319, 20046, 24999, 25436, 25011, 24013, 23172, 22995, 22937, 22978, 
    23255, 23872, 24881, 26141, 27005, 23174, 26327, 26375, 25903, 25440, 
    24871, 24274,
  20047, 19654, 25251, 25492, 24959, 23934, 23146, 22981, 22978, 22948, 
    23270, 23845, 24995, 26238, 27337, 23515, 26386, 26285, 25800, 25348, 
    24795, 24222,
  28064, 28015, 28007, 27271, 25892, 24208, 22712, 22299, 22212, 22526, 
    22973, 23674, 24687, 25683, 26806, 28649, 29009, 28065, 27315, 26544, 
    25600, 24513,
  28062, 28034, 28004, 27349, 26028, 24327, 22812, 22296, 22159, 22545, 
    22917, 23606, 24572, 25766, 26466, 28600, 28999, 28040, 27412, 26593, 
    25511, 24385,
  28057, 28088, 28022, 27359, 26139, 24422, 22876, 22364, 22198, 22473, 
    22903, 23622, 24730, 25880, 26487, 28554, 29029, 28029, 27303, 26537, 
    25513, 24426,
  28015, 28113, 27979, 27374, 26195, 24504, 22974, 22379, 22181, 22568, 
    22882, 23609, 24535, 25899, 26681, 28503, 28924, 27897, 27175, 26388, 
    25404, 24265,
  27999, 28127, 27910, 27467, 26263, 24636, 23049, 22442, 22213, 22519, 
    22950, 23545, 24536, 25810, 26599, 28371, 28687, 27735, 26941, 26226, 
    25164, 24151,
  27954, 28089, 27872, 27397, 26293, 24686, 23089, 22459, 22201, 22471, 
    22933, 23573, 24500, 25760, 26725, 28262, 28660, 27673, 26867, 26034, 
    25029, 24110,
  27869, 27979, 27766, 27368, 26401, 24796, 23161, 22507, 22247, 22514, 
    22923, 23435, 24447, 25689, 26669, 28218, 28604, 27704, 26928, 26115, 
    25107, 24117,
  27764, 27843, 27757, 27397, 26443, 24818, 23227, 22564, 22259, 22492, 
    22926, 23458, 24467, 25779, 27054, 28172, 28597, 27603, 26905, 26157, 
    25094, 24150,
  27654, 27722, 27654, 27350, 26468, 24901, 23265, 22583, 22268, 22515, 
    22793, 23481, 24486, 25777, 26366, 28099, 28472, 27375, 26674, 26015, 
    25075, 24157,
  27536, 27625, 27562, 27287, 26472, 24962, 23336, 22642, 22254, 22454, 
    22890, 23488, 24310, 25548, 26579, 27949, 28275, 27241, 26500, 25854, 
    24999, 24265,
  27416, 27523, 27423, 27233, 26441, 24995, 23407, 22623, 22302, 22542, 
    22911, 23401, 24340, 25584, 26626, 27809, 28013, 26938, 26249, 25580, 
    24991, 24243,
  27322, 27416, 27286, 27140, 26435, 25017, 23432, 22671, 22341, 22522, 
    22915, 23451, 24460, 25595, 26713, 27639, 27785, 26632, 25937, 25409, 
    24792, 24142,
  27267, 27333, 27172, 27049, 26374, 25026, 23455, 22693, 22282, 22508, 
    22910, 23472, 24302, 25657, 26797, 27401, 27448, 26359, 25753, 25220, 
    24555, 23993,
  27264, 27302, 27051, 26913, 26315, 25018, 23555, 22726, 22354, 22479, 
    22915, 23376, 24444, 25490, 26769, 27192, 27108, 26253, 25724, 25186, 
    24540, 23910,
  27273, 27323, 26942, 26854, 26250, 25028, 23561, 22764, 22412, 22506, 
    22837, 23471, 24342, 25715, 26959, 26832, 26453, 26035, 25576, 25115, 
    24467, 23940,
  27619, 27567, 27082, 26816, 26213, 25002, 23583, 22707, 22293, 22394, 
    22784, 23403, 24430, 25486, 26732, 26735, 25572, 25563, 25298, 24933, 
    24299, 23806,
  27536, 27489, 27081, 26899, 26229, 25083, 23604, 22760, 22334, 22491, 
    22827, 23342, 24202, 25383, 26795, 26885, 25801, 25628, 25401, 25001, 
    24439, 23940,
  27058, 27118, 27044, 26931, 26421, 25204, 23689, 22837, 22436, 22440, 
    22917, 23369, 24286, 25471, 26522, 27106, 26874, 26228, 25690, 25197, 
    24595, 24027,
  26943, 26980, 26881, 26896, 26446, 25260, 23699, 22890, 22424, 22420, 
    22982, 23470, 24426, 25616, 26520, 27185, 27287, 26422, 25800, 25221, 
    24626, 23993,
  26881, 26894, 26650, 26722, 26401, 25307, 23789, 22901, 22446, 22532, 
    22811, 23387, 24264, 25424, 26546, 27023, 27243, 26366, 25779, 25145, 
    24504, 23953,
  26881, 26880, 26799, 26817, 26433, 25260, 23776, 22988, 22464, 22460, 
    22841, 23390, 24230, 25556, 26768, 27146, 27294, 26322, 25712, 25060, 
    24448, 23866,
  26922, 26915, 26978, 26944, 26500, 25320, 23796, 22997, 22512, 22484, 
    22902, 23383, 24279, 25340, 26778, 27379, 27265, 26241, 25601, 25104, 
    24492, 23872,
  26959, 26960, 26944, 26853, 26494, 25315, 23817, 23001, 22499, 22513, 
    22729, 23309, 24275, 25446, 26296, 27414, 27175, 26257, 25637, 25041, 
    24409, 23824,
  26975, 26996, 26810, 26850, 26434, 25320, 23818, 23000, 22540, 22537, 
    22810, 23338, 24248, 25470, 26809, 27318, 27200, 26281, 25701, 25064, 
    24420, 23950,
  27003, 27026, 26874, 26870, 26430, 25309, 23871, 23051, 22534, 22446, 
    22876, 23360, 24234, 25424, 26689, 27316, 27157, 26350, 25713, 25201, 
    24571, 23887,
  27062, 27085, 27006, 26887, 26446, 25307, 23845, 23062, 22518, 22528, 
    22868, 23279, 24202, 25465, 26356, 27354, 27104, 26232, 25741, 25255, 
    24588, 23852,
  27127, 27172, 26940, 26913, 26429, 25366, 23908, 23052, 22589, 22533, 
    22918, 23357, 24249, 25446, 26657, 27306, 27019, 26210, 25704, 25178, 
    24485, 23951,
  27158, 27257, 26865, 26765, 26357, 25347, 23890, 23065, 22609, 22527, 
    22850, 23427, 24271, 25312, 26453, 27101, 26969, 26239, 25803, 25256, 
    24656, 23850,
  27139, 27282, 26849, 26744, 26326, 25333, 23922, 23123, 22592, 22561, 
    22900, 23395, 24300, 25353, 26261, 27064, 26865, 26326, 25827, 25255, 
    24565, 24004,
  27076, 27216, 26849, 26739, 26328, 25342, 23939, 23120, 22631, 22549, 
    22766, 23398, 24246, 25288, 26645, 27035, 26912, 26316, 25874, 25304, 
    24603, 24017,
  26947, 27046, 26779, 26719, 26281, 25329, 23947, 23102, 22599, 22512, 
    22753, 23315, 24175, 25344, 26621, 27025, 26853, 26240, 25746, 25221, 
    24609, 23952,
  26707, 26778, 26765, 26665, 26296, 25348, 23990, 23169, 22637, 22532, 
    22803, 23375, 24267, 25406, 26645, 26988, 26941, 26272, 25855, 25315, 
    24648, 24039,
  26322, 26407, 26642, 26590, 26257, 25300, 23970, 23185, 22642, 22563, 
    22807, 23344, 24397, 25352, 26513, 26982, 26923, 26349, 25820, 25251, 
    24655, 24085,
  25840, 25947, 26529, 26542, 26238, 25311, 24015, 23182, 22685, 22562, 
    22895, 23317, 24231, 25458, 26665, 26888, 26904, 26363, 25888, 25315, 
    24673, 24139,
  25362, 25478, 26335, 26434, 26170, 25327, 24007, 23232, 22644, 22578, 
    22827, 23307, 24207, 25434, 26528, 26748, 26813, 26222, 25776, 25172, 
    24602, 24004,
  24992, 25104, 26181, 26322, 26187, 25295, 24015, 23200, 22658, 22611, 
    22919, 23422, 24183, 25340, 26334, 26623, 26565, 26034, 25584, 25149, 
    24615, 23984,
  24802, 24901, 25999, 26230, 26106, 25319, 24052, 23231, 22689, 22630, 
    22887, 23432, 24084, 25585, 26682, 26435, 26240, 25772, 25425, 24985, 
    24462, 24020,
  25127, 25042, 26226, 26370, 26148, 25291, 24014, 23124, 22614, 22633, 
    22820, 23275, 24214, 25318, 26450, 26476, 25879, 25429, 25183, 24829, 
    24351, 23901,
  25230, 25080, 26184, 26324, 26114, 25310, 24000, 23156, 22614, 22616, 
    22868, 23374, 24229, 25376, 26268, 26399, 25918, 25444, 25155, 24785, 
    24364, 23914,
  24979, 24916, 25854, 26090, 26101, 25349, 24073, 23216, 22779, 22605, 
    22865, 23411, 24207, 25465, 26218, 26145, 26051, 25524, 25168, 24798, 
    24418, 23782,
  24909, 24844, 25841, 26113, 26097, 25336, 24054, 23249, 22735, 22608, 
    22849, 23346, 24119, 25422, 26306, 26114, 26237, 25667, 25327, 24885, 
    24521, 24031,
  24673, 24628, 25756, 26069, 26061, 25300, 24070, 23226, 22746, 22619, 
    22861, 23320, 24162, 25386, 26419, 25999, 26315, 25862, 25464, 24990, 
    24496, 24046,
  24344, 24314, 25601, 25961, 25983, 25282, 24062, 23260, 22706, 22616, 
    22915, 23360, 24245, 25333, 26606, 25760, 25825, 25719, 25408, 25123, 
    24572, 24020,
  24052, 24009, 25348, 25790, 25903, 25304, 24051, 23284, 22774, 22642, 
    22912, 23331, 24439, 25393, 26321, 25402, 25223, 25385, 25259, 25048, 
    24605, 24040,
  24196, 23995, 25491, 25896, 25904, 25243, 24055, 23171, 22707, 22595, 
    22828, 23363, 24157, 25238, 26478, 25377, 25114, 25154, 25099, 24809, 
    24433, 23974,
  24183, 23975, 25512, 25976, 25897, 25221, 24014, 23177, 22681, 22586, 
    22802, 23317, 24067, 25248, 26629, 25377, 25319, 25284, 25244, 24940, 
    24452, 24068,
  23988, 23926, 25404, 25835, 25989, 25312, 24042, 23251, 22740, 22567, 
    22904, 23375, 24251, 25367, 26753, 25262, 25666, 25497, 25350, 25076, 
    24528, 24131,
  24433, 24254, 25714, 26060, 26014, 25282, 24007, 23189, 22701, 22603, 
    22862, 23416, 24045, 25175, 26406, 25519, 25681, 25508, 25348, 24990, 
    24459, 24041,
  24600, 24435, 25684, 26017, 25988, 25254, 24058, 23162, 22669, 22661, 
    22888, 23305, 24018, 25227, 26488, 25457, 25662, 25494, 25320, 24978, 
    24580, 24081,
  24742, 24582, 25862, 26095, 25994, 25277, 24021, 23203, 22689, 22641, 
    22911, 23289, 24070, 25380, 26469, 25580, 25681, 25552, 25328, 25021, 
    24478, 24041,
  24517, 24499, 25596, 25999, 25983, 25336, 24077, 23288, 22790, 22725, 
    22950, 23375, 24217, 25348, 26566, 25461, 26070, 25726, 25460, 25179, 
    24608, 24094,
  24457, 24459, 25525, 25959, 26020, 25348, 24044, 23285, 22809, 22668, 
    23004, 23426, 24137, 25352, 26554, 25484, 26200, 25831, 25458, 25052, 
    24626, 24109,
  24536, 24444, 25748, 26095, 26022, 25268, 24014, 23159, 22721, 22712, 
    22990, 23383, 24208, 25444, 26285, 25644, 26329, 25862, 25466, 24959, 
    24497, 24021,
  23857, 23954, 25304, 25830, 25975, 25285, 24028, 23284, 22819, 22726, 
    22997, 23401, 24313, 25425, 26415, 25183, 26601, 26131, 25629, 25199, 
    24532, 24116,
  23343, 23491, 24842, 25578, 25845, 25298, 24039, 23284, 22807, 22760, 
    23014, 23416, 24221, 25454, 26610, 24568, 26291, 26290, 25774, 25199, 
    24672, 24190,
  22752, 22939, 24590, 25408, 25782, 25244, 24027, 23293, 22846, 22721, 
    22967, 23474, 24221, 25452, 26366, 24217, 26241, 26394, 25825, 25305, 
    24672, 24210,
  22109, 22310, 24579, 25387, 25799, 25234, 24049, 23304, 22848, 22791, 
    22856, 23403, 24261, 25457, 26472, 24372, 26582, 26538, 25935, 25332, 
    24724, 24216,
  21403, 21574, 24295, 25196, 25690, 25232, 24037, 23256, 22810, 22668, 
    23074, 23418, 24307, 25443, 27025, 24106, 26486, 26629, 26004, 25443, 
    24755, 24144,
  20622, 20757, 23891, 24951, 25618, 25195, 24003, 23277, 22846, 22756, 
    23045, 23404, 24285, 25320, 26499, 23679, 26159, 26664, 26107, 25443, 
    24762, 24198,
  19828, 19937, 23590, 24737, 25525, 25164, 23942, 23257, 22856, 22769, 
    23019, 23423, 24320, 25487, 26532, 23635, 26391, 26769, 26188, 25625, 
    24821, 24278,
  19173, 19267, 22932, 24380, 25364, 25099, 23953, 23252, 22842, 22744, 
    23013, 23368, 24258, 25654, 26343, 23074, 26200, 26753, 26303, 25636, 
    25015, 24340,
  18765, 18860, 22378, 24017, 25220, 25067, 23988, 23261, 22833, 22768, 
    23023, 23423, 24359, 25550, 26651, 22404, 25661, 26742, 26298, 25719, 
    24926, 24414,
  18621, 18730, 22054, 23826, 25107, 25026, 23912, 23262, 22809, 22764, 
    22946, 23321, 24198, 25553, 26549, 22165, 25294, 26741, 26334, 25789, 
    25011, 24284,
  18683, 18810, 22080, 23796, 25047, 24986, 23923, 23218, 22882, 22795, 
    22974, 23458, 24258, 25513, 26345, 22062, 24962, 26716, 26355, 25826, 
    25025, 24454,
  18869, 19041, 22073, 23773, 25017, 24921, 23907, 23263, 22845, 22787, 
    23022, 23466, 24220, 25268, 26602, 22020, 24801, 26579, 26382, 25807, 
    25095, 24474,
  19134, 19370, 22188, 23828, 25013, 24935, 23893, 23232, 22878, 22821, 
    23025, 23414, 24311, 25480, 26672, 22148, 24938, 26672, 26399, 25906, 
    25178, 24554,
  19448, 19735, 22494, 24029, 25129, 24933, 23857, 23214, 22842, 22812, 
    23102, 23370, 24485, 25411, 26492, 22372, 25167, 26708, 26513, 25979, 
    25211, 24675,
  19716, 20026, 22931, 24300, 25206, 24926, 23878, 23197, 22873, 22820, 
    23107, 23458, 24312, 25522, 26696, 22752, 25403, 26704, 26493, 26026, 
    25236, 24544,
  19807, 20125, 23270, 24476, 25297, 24921, 23818, 23213, 22821, 22789, 
    23053, 23572, 24345, 25644, 26484, 23086, 25618, 26741, 26492, 26079, 
    25339, 24679,
  19634, 19962, 23381, 24551, 25285, 24915, 23849, 23214, 22891, 22826, 
    23065, 23591, 24271, 25423, 26673, 23224, 25736, 26744, 26454, 25927, 
    25290, 24687,
  19210, 19559, 23213, 24487, 25242, 24830, 23793, 23192, 22857, 22805, 
    23050, 23496, 24458, 25556, 26721, 23029, 25663, 26656, 26449, 25904, 
    25287, 24540,
  18665, 19011, 22882, 24332, 25176, 24871, 23796, 23170, 22854, 22859, 
    23089, 23490, 24382, 25791, 26671, 22672, 25519, 26668, 26429, 25939, 
    25331, 24679,
  18126, 18444, 22383, 24041, 25106, 24817, 23773, 23215, 22888, 22822, 
    23076, 23511, 24424, 25641, 26493, 22118, 25336, 26659, 26400, 26008, 
    25385, 24741,
  17661, 17944, 22019, 23809, 25024, 24750, 23741, 23170, 22892, 22861, 
    22934, 23465, 24354, 25465, 26771, 21542, 24830, 26584, 26412, 25875, 
    25341, 24587,
  17249, 17536, 21811, 23731, 25000, 24748, 23748, 23195, 22900, 22853, 
    23114, 23633, 24442, 25684, 26895, 21293, 24696, 26603, 26316, 25903, 
    25261, 24582,
  16868, 17166, 21698, 23724, 24999, 24782, 23724, 23201, 22924, 22921, 
    23081, 23565, 24434, 25713, 26943, 21135, 24803, 26651, 26351, 25860, 
    25254, 24785,
  16503, 16807, 21643, 23694, 24979, 24689, 23687, 23177, 22940, 22909, 
    23229, 23623, 24420, 25576, 26569, 21147, 24960, 26613, 26268, 25819, 
    25192, 24723,
  16210, 16477, 21692, 23742, 25029, 24662, 23687, 23132, 22932, 22911, 
    23141, 23498, 24544, 25626, 26593, 21155, 25104, 26632, 26272, 25734, 
    25238, 24524,
  16027, 16252, 21847, 23777, 25036, 24658, 23654, 23172, 22917, 22884, 
    23154, 23539, 24502, 25807, 26880, 21234, 25210, 26593, 26220, 25793, 
    25215, 24626,
  16027, 16209, 21946, 23851, 25000, 24619, 23611, 23162, 22951, 22919, 
    23147, 23559, 24490, 25588, 27009, 21335, 25213, 26638, 26290, 25862, 
    25286, 24727,
  16269, 16473, 22074, 23956, 25047, 24617, 23603, 23117, 22943, 22882, 
    23105, 23622, 24579, 25865, 27072, 21462, 25414, 26637, 26300, 25871, 
    25320, 24748,
  16889, 17115, 22390, 24170, 25068, 24612, 23609, 23132, 22934, 22923, 
    23165, 23637, 24617, 25818, 26913, 21625, 25465, 26618, 26267, 25805, 
    25187, 24656,
  17929, 18137, 22914, 24454, 25171, 24602, 23572, 23155, 22991, 22949, 
    23087, 23678, 24612, 26044, 27270, 22026, 25523, 26549, 26179, 25706, 
    25086, 24537,
  19246, 19371, 23796, 24892, 25240, 24555, 23532, 23121, 22958, 22983, 
    23201, 23656, 24591, 25925, 27150, 22943, 25801, 26605, 26193, 25724, 
    25093, 24464,
  20510, 20559, 24521, 25237, 25326, 24543, 23530, 23117, 22989, 22989, 
    23228, 23641, 24664, 25848, 26971, 23823, 26144, 26573, 26187, 25743, 
    25079, 24553,
  21474, 21488, 24755, 25373, 25356, 24498, 23548, 23062, 23023, 23006, 
    23096, 23684, 24582, 25975, 26779, 24157, 26121, 26551, 26151, 25650, 
    25024, 24474,
  22101, 22142, 24626, 25300, 25300, 24421, 23492, 23108, 22989, 22996, 
    23273, 23624, 24619, 26074, 26893, 23896, 26110, 26501, 26128, 25586, 
    25049, 24481,
  22558, 22650, 24616, 25346, 25297, 24364, 23437, 23087, 22967, 23009, 
    23345, 23672, 24562, 26214, 27307, 23716, 25994, 26501, 26100, 25747, 
    25172, 24688,
  22985, 23104, 25074, 25606, 25321, 24344, 23442, 23067, 22944, 22979, 
    23243, 23825, 24698, 26006, 27066, 24230, 26434, 26519, 26068, 25716, 
    25108, 24535,
  23309, 23433, 25605, 25785, 25369, 24387, 23389, 23090, 22993, 23060, 
    23247, 23850, 24731, 26029, 27130, 24882, 26622, 26566, 26131, 25655, 
    25090, 24562,
  23325, 23451, 25676, 25810, 25325, 24232, 23370, 23076, 22937, 23023, 
    23175, 23773, 24758, 26123, 26956, 25236, 26625, 26515, 26135, 25720, 
    25029, 24403,
  22941, 23081, 25633, 25763, 25226, 24208, 23303, 23046, 22983, 23019, 
    23222, 23742, 24818, 26263, 27128, 25254, 26614, 26473, 26050, 25545, 
    24942, 24318,
  22237, 22340, 25362, 25622, 25147, 24160, 23253, 23042, 22990, 22986, 
    23282, 23852, 24876, 26304, 27106, 24686, 26632, 26416, 25971, 25497, 
    24880, 24287,
  21420, 21361, 24989, 25445, 25077, 24090, 23231, 22993, 22985, 23011, 
    23222, 23789, 24822, 26381, 26981, 23475, 26422, 26363, 25944, 25526, 
    24864, 24351,
  20683, 20418, 24990, 25420, 25000, 24034, 23200, 23015, 22971, 23025, 
    23331, 23892, 24923, 26416, 26846, 23170, 26333, 26315, 25872, 25491, 
    24835, 24308,
  20391, 20011, 25209, 25480, 24953, 23951, 23171, 23013, 22954, 23024, 
    23272, 23850, 24985, 26368, 27112, 23579, 26428, 26247, 25747, 25250, 
    24645, 24056,
  28031, 27977, 27974, 27308, 25909, 24172, 22762, 22277, 22182, 22555, 
    22902, 23701, 24665, 25774, 26841, 28685, 29138, 28071, 27403, 26648, 
    25518, 24486,
  28035, 28002, 27979, 27381, 26037, 24316, 22817, 22344, 22202, 22465, 
    22998, 23611, 24537, 25785, 26734, 28622, 29073, 28061, 27354, 26561, 
    25531, 24512,
  28044, 28065, 27949, 27388, 26128, 24380, 22883, 22355, 22197, 22493, 
    22992, 23577, 24680, 25890, 26885, 28571, 28978, 27970, 27288, 26562, 
    25456, 24386,
  28011, 28092, 27951, 27395, 26200, 24529, 23018, 22394, 22198, 22500, 
    22901, 23535, 24598, 25560, 26535, 28542, 28873, 27874, 27132, 26399, 
    25342, 24312,
  27993, 28101, 27874, 27424, 26255, 24594, 23048, 22413, 22195, 22511, 
    22862, 23612, 24473, 25828, 26734, 28413, 28723, 27800, 27063, 26269, 
    25139, 24298,
  27940, 28056, 27787, 27360, 26278, 24726, 23130, 22489, 22232, 22493, 
    22894, 23585, 24615, 25648, 26576, 28290, 28659, 27672, 26899, 26119, 
    25062, 24124,
  27839, 27936, 27694, 27429, 26331, 24745, 23165, 22502, 22238, 22485, 
    22896, 23457, 24448, 25754, 26576, 28221, 28529, 27588, 26774, 26119, 
    25050, 24137,
  27704, 27775, 27649, 27356, 26429, 24827, 23247, 22585, 22249, 22489, 
    22864, 23460, 24461, 25620, 26693, 28183, 28402, 27363, 26565, 25828, 
    24949, 24003,
  27552, 27611, 27561, 27322, 26426, 24879, 23302, 22592, 22257, 22474, 
    22873, 23443, 24364, 25577, 26741, 28063, 28297, 27094, 26390, 25734, 
    24822, 24096,
  27391, 27464, 27435, 27222, 26400, 24912, 23307, 22628, 22318, 22491, 
    22810, 23566, 24408, 25565, 26871, 27869, 28049, 26937, 26291, 25561, 
    24930, 24117,
  27251, 27334, 27210, 27048, 26353, 24920, 23375, 22657, 22339, 22543, 
    22792, 23525, 24234, 25705, 26710, 27596, 27657, 26578, 25965, 25448, 
    24731, 24109,
  27169, 27235, 27066, 26868, 26284, 24968, 23465, 22695, 22372, 22493, 
    22879, 23461, 24447, 25709, 26903, 27217, 27254, 26292, 25722, 25190, 
    24609, 23848,
  27152, 27187, 26963, 26812, 26243, 24926, 23477, 22737, 22322, 22453, 
    22862, 23436, 24464, 25464, 26416, 26976, 26395, 25969, 25518, 25100, 
    24499, 23940,
  27192, 27194, 26940, 26821, 26218, 25015, 23523, 22768, 22376, 22532, 
    22925, 23525, 24318, 25506, 26444, 26826, 26429, 25965, 25563, 25122, 
    24459, 23985,
  27227, 27238, 26871, 26764, 26271, 25017, 23521, 22809, 22426, 22468, 
    22878, 23487, 24489, 25581, 26644, 26712, 26128, 25912, 25588, 25102, 
    24519, 23933,
  27573, 27485, 27053, 26749, 26165, 25014, 23551, 22740, 22313, 22397, 
    22825, 23388, 24293, 25162, 26510, 26710, 25484, 25433, 25289, 24876, 
    24371, 23720,
  27475, 27400, 27124, 26818, 26245, 25098, 23603, 22716, 22351, 22448, 
    22828, 23420, 24187, 25616, 26229, 26828, 25484, 25368, 25282, 25006, 
    24440, 23967,
  26982, 27027, 26907, 26885, 26396, 25218, 23681, 22853, 22418, 22500, 
    22816, 23460, 24211, 25259, 26878, 27020, 26667, 26076, 25674, 25221, 
    24621, 23941,
  26863, 26900, 26715, 26794, 26356, 25193, 23711, 22844, 22456, 22518, 
    22832, 23389, 24218, 25315, 26541, 27070, 27317, 26372, 25860, 25145, 
    24627, 24073,
  26806, 26831, 26587, 26712, 26361, 25209, 23725, 22923, 22501, 22499, 
    22869, 23371, 24283, 25492, 26675, 26939, 27335, 26380, 25729, 25113, 
    24512, 23947,
  26807, 26831, 26782, 26772, 26387, 25232, 23778, 22995, 22527, 22535, 
    22860, 23401, 24281, 25442, 26416, 27166, 27237, 26250, 25654, 25146, 
    24456, 23879,
  26840, 26870, 26925, 26874, 26368, 25267, 23781, 22989, 22491, 22511, 
    22729, 23334, 24152, 25268, 26782, 27309, 26976, 26126, 25619, 25097, 
    24481, 23846,
  26873, 26917, 26876, 26780, 26388, 25273, 23833, 22961, 22512, 22499, 
    22832, 23441, 24387, 25385, 26768, 27335, 26768, 26026, 25581, 25039, 
    24474, 23884,
  26910, 26958, 26768, 26767, 26353, 25348, 23831, 23007, 22522, 22592, 
    22912, 23459, 24229, 25323, 26451, 27273, 26721, 26043, 25638, 25193, 
    24504, 23917,
  26977, 26995, 26847, 26806, 26376, 25292, 23836, 23028, 22545, 22460, 
    22849, 23349, 24255, 25519, 26246, 27324, 26894, 26206, 25725, 25231, 
    24579, 23934,
  27064, 27058, 26953, 26938, 26432, 25326, 23882, 23080, 22586, 22496, 
    22865, 23421, 24295, 25296, 26559, 27441, 27171, 26434, 25891, 25359, 
    24627, 23966,
  27130, 27143, 26917, 26888, 26416, 25328, 23903, 23070, 22545, 22508, 
    22817, 23336, 24175, 25342, 26467, 27353, 27229, 26449, 25929, 25251, 
    24632, 23978,
  27140, 27220, 26868, 26822, 26340, 25283, 23934, 23115, 22597, 22536, 
    22910, 23395, 24168, 25326, 26743, 27222, 27024, 26477, 25912, 25361, 
    24637, 24031,
  27097, 27232, 26831, 26760, 26310, 25298, 23914, 23118, 22593, 22582, 
    22770, 23288, 24165, 25400, 26723, 27158, 26975, 26371, 25943, 25366, 
    24655, 24131,
  27010, 27150, 26804, 26715, 26306, 25318, 23906, 23118, 22610, 22567, 
    22915, 23370, 24292, 25325, 26489, 27050, 27047, 26569, 25941, 25340, 
    24700, 24245,
  26854, 26962, 26803, 26695, 26293, 25282, 23945, 23144, 22625, 22576, 
    22939, 23286, 24211, 25510, 26768, 27038, 26971, 26456, 25985, 25437, 
    24738, 24025,
  26584, 26672, 26756, 26724, 26267, 25312, 23953, 23143, 22616, 22515, 
    22875, 23337, 24234, 25418, 26320, 27038, 26989, 26453, 26019, 25394, 
    24706, 24099,
  26174, 26272, 26657, 26631, 26254, 25300, 23983, 23165, 22688, 22572, 
    22860, 23307, 24125, 25228, 26744, 26957, 26929, 26443, 26046, 25399, 
    24719, 24152,
  25673, 25784, 26351, 26491, 26144, 25286, 24017, 23168, 22648, 22571, 
    22851, 23382, 24074, 25419, 26276, 26846, 26816, 26406, 25982, 25494, 
    24789, 24145,
  25174, 25297, 26243, 26357, 26104, 25282, 24009, 23141, 22658, 22584, 
    22908, 23287, 24402, 25393, 26540, 26778, 26793, 26425, 26010, 25488, 
    24769, 24247,
  24771, 24915, 26118, 26220, 26075, 25315, 24020, 23200, 22730, 22685, 
    22866, 23358, 24249, 25396, 26601, 26622, 26601, 26206, 25760, 25327, 
    24724, 24145,
  24869, 24893, 26226, 26373, 26049, 25246, 24020, 23116, 22654, 22532, 
    22775, 23292, 24134, 25313, 26415, 26671, 26185, 25625, 25416, 24996, 
    24531, 24022,
  24518, 24643, 25825, 26064, 26047, 25289, 24026, 23221, 22735, 22613, 
    22886, 23343, 24222, 25339, 26357, 26187, 25794, 25396, 25195, 24866, 
    24469, 23967,
  24635, 24677, 25717, 26047, 26037, 25307, 24038, 23224, 22740, 22684, 
    22885, 23344, 24209, 25378, 26487, 25968, 25546, 25297, 25099, 24834, 
    24354, 23895,
  24760, 24723, 25710, 26042, 26029, 25316, 24044, 23252, 22700, 22640, 
    22954, 23362, 24176, 25311, 26854, 25889, 25696, 25459, 25229, 24902, 
    24393, 23843,
  24761, 24699, 25729, 26066, 26083, 25354, 24036, 23287, 22752, 22654, 
    22836, 23381, 24151, 25264, 26344, 25907, 26087, 25782, 25505, 25095, 
    24565, 24004,
  24599, 24547, 25616, 25991, 26007, 25326, 24026, 23266, 22757, 22617, 
    22899, 23236, 24178, 25246, 26826, 25899, 26538, 26063, 25669, 25169, 
    24554, 23966,
  24332, 24297, 25475, 25927, 26075, 25333, 24068, 23272, 22825, 22691, 
    22926, 23377, 24213, 25547, 26201, 25732, 26466, 26016, 25566, 25072, 
    24631, 24034,
  24084, 24049, 25436, 25913, 25995, 25361, 24070, 23265, 22771, 22625, 
    22962, 23337, 24126, 25421, 26415, 25537, 26312, 25912, 25596, 25165, 
    24600, 24134,
  23941, 23907, 25282, 25810, 26004, 25296, 24080, 23269, 22762, 22629, 
    22860, 23287, 24195, 25296, 26328, 25314, 26201, 25897, 25546, 25159, 
    24650, 24093,
  24235, 24072, 25517, 25901, 25985, 25252, 24019, 23159, 22671, 22610, 
    22895, 23360, 24156, 25337, 26422, 25399, 26091, 25776, 25498, 25094, 
    24612, 24068,
  24318, 24168, 25606, 25944, 25974, 25316, 24047, 23204, 22715, 22649, 
    22854, 23317, 24094, 25472, 26613, 25471, 25997, 25710, 25367, 25020, 
    24562, 24021,
  24450, 24308, 25689, 25995, 26016, 25280, 24057, 23219, 22703, 22655, 
    22829, 23278, 24013, 25472, 26610, 25527, 25848, 25573, 25367, 25063, 
    24441, 24075,
  24593, 24460, 25798, 26022, 26001, 25305, 24019, 23213, 22727, 22624, 
    22900, 23319, 24047, 25376, 26194, 25571, 25804, 25479, 25325, 24957, 
    24492, 24115,
  24435, 24446, 25607, 25959, 26041, 25336, 24071, 23266, 22848, 22691, 
    22979, 23369, 24280, 25276, 26787, 25543, 26143, 25826, 25462, 25045, 
    24597, 24061,
  24499, 24539, 25697, 26010, 26066, 25342, 24051, 23263, 22809, 22616, 
    22962, 23372, 24312, 25500, 26484, 25676, 26150, 25857, 25444, 25116, 
    24565, 24020,
  24776, 24715, 25862, 26149, 26037, 25266, 24009, 23189, 22741, 22644, 
    22909, 23327, 24131, 25306, 26662, 25689, 26110, 25776, 25381, 24989, 
    24460, 24121,
  24641, 24617, 25837, 26041, 25997, 25246, 24005, 23162, 22735, 22652, 
    22900, 23296, 24220, 25418, 26572, 25591, 26159, 25782, 25374, 25032, 
    24485, 24055,
  24080, 24228, 25523, 25886, 25999, 25266, 24023, 23284, 22815, 22695, 
    22938, 23299, 24276, 25426, 26337, 25418, 26469, 26153, 25682, 25135, 
    24629, 24082,
  23684, 23865, 25461, 25912, 25983, 25236, 24058, 23320, 22792, 22691, 
    22944, 23377, 23983, 25349, 26443, 25319, 26675, 26369, 25820, 25266, 
    24641, 24103,
  23149, 23365, 25196, 25724, 25876, 25283, 24040, 23268, 22848, 22692, 
    22877, 23420, 24161, 25497, 26712, 24964, 26613, 26503, 25900, 25310, 
    24591, 24149,
  22444, 22682, 24832, 25499, 25838, 25276, 24003, 23259, 22835, 22691, 
    22925, 23334, 24163, 25457, 26450, 24719, 26569, 26588, 25974, 25387, 
    24718, 24203,
  21525, 21753, 24412, 25256, 25731, 25255, 24014, 23265, 22828, 22725, 
    23018, 23405, 24351, 25490, 26599, 24314, 26441, 26644, 26057, 25443, 
    24667, 24157,
  20390, 20612, 23645, 24874, 25586, 25142, 23985, 23301, 22816, 22651, 
    22946, 23325, 24420, 25404, 26295, 23721, 26384, 26757, 26154, 25616, 
    24847, 24238,
  19151, 19377, 22744, 24231, 25281, 25043, 23975, 23272, 22846, 22732, 
    22974, 23376, 24176, 25468, 26745, 22755, 25903, 26740, 26271, 25699, 
    24880, 24271,
  18045, 18273, 21934, 23778, 25095, 25010, 23938, 23229, 22836, 22772, 
    22988, 23399, 24210, 25350, 26509, 21868, 25376, 26766, 26301, 25759, 
    24887, 24171,
  17277, 17500, 21675, 23539, 24999, 25014, 23942, 23253, 22826, 22743, 
    23010, 23435, 24245, 25610, 26487, 21543, 25405, 26742, 26324, 25712, 
    24959, 24354,
  16944, 17151, 21651, 23558, 24987, 24935, 23936, 23248, 22829, 22761, 
    22932, 23367, 24118, 25455, 26891, 21529, 25237, 26689, 26422, 25850, 
    25139, 24345,
  17016, 17204, 21794, 23565, 24981, 24910, 23929, 23248, 22835, 22777, 
    23010, 23359, 24301, 25540, 26596, 21519, 25180, 26701, 26429, 25937, 
    25146, 24487,
  17391, 17583, 21812, 23561, 24974, 24959, 23902, 23264, 22835, 22796, 
    22932, 23470, 24370, 25608, 26446, 21563, 25037, 26716, 26450, 25992, 
    25204, 24467,
  17962, 18184, 22002, 23714, 24984, 24871, 23867, 23195, 22895, 22841, 
    23018, 23475, 24283, 25370, 26394, 21768, 25068, 26772, 26446, 26029, 
    25235, 24581,
  18631, 18879, 22484, 23987, 25069, 24905, 23845, 23191, 22903, 22762, 
    22920, 23422, 24097, 25253, 26732, 22230, 25210, 26736, 26491, 26022, 
    25301, 24460,
  19254, 19518, 23042, 24314, 25174, 24881, 23851, 23204, 22855, 22746, 
    22991, 23412, 24256, 25518, 26264, 22872, 25583, 26739, 26450, 26018, 
    25307, 24664,
  19675, 19960, 23404, 24552, 25266, 24885, 23842, 23196, 22873, 22821, 
    22980, 23447, 24167, 25319, 26679, 23342, 25772, 26625, 26455, 25947, 
    25372, 24638,
  19794, 20122, 23530, 24601, 25308, 24898, 23785, 23209, 22846, 22835, 
    23029, 23421, 24300, 25491, 26728, 23455, 25810, 26759, 26439, 26006, 
    25284, 24646,
  19605, 19995, 23375, 24577, 25276, 24861, 23793, 23204, 22888, 22819, 
    23037, 23500, 24411, 25738, 26948, 23251, 25626, 26763, 26522, 26015, 
    25358, 24755,
  19203, 19625, 23041, 24365, 25247, 24857, 23759, 23191, 22898, 22853, 
    23010, 23392, 24280, 25438, 26650, 22891, 25412, 26668, 26454, 25906, 
    25345, 24718,
  18703, 19102, 22737, 24181, 25118, 24817, 23760, 23211, 22896, 22880, 
    23076, 23650, 24394, 25646, 26505, 22462, 25298, 26666, 26460, 25938, 
    25353, 24787,
  18186, 18524, 22389, 23993, 25073, 24785, 23723, 23176, 22910, 22896, 
    22975, 23477, 24407, 25559, 26870, 21945, 25022, 26656, 26348, 25850, 
    25266, 24660,
  17664, 17972, 22135, 23920, 25041, 24760, 23719, 23196, 22879, 22854, 
    23041, 23562, 24441, 25625, 26674, 21671, 25064, 26588, 26308, 25846, 
    25204, 24648,
  17148, 17451, 21931, 23751, 25018, 24732, 23729, 23203, 22888, 22871, 
    23151, 23587, 24394, 25651, 26719, 21387, 24914, 26615, 26294, 25778, 
    25287, 24651,
  16638, 16954, 21764, 23709, 24965, 24639, 23646, 23149, 22898, 22898, 
    23096, 23506, 24456, 25520, 26709, 21218, 24891, 26599, 26232, 25781, 
    25244, 24649,
  16205, 16492, 21692, 23691, 24977, 24653, 23668, 23168, 22951, 22902, 
    23065, 23460, 24385, 25624, 26675, 21168, 25128, 26603, 26298, 25788, 
    25207, 24664,
  15913, 16158, 21818, 23816, 25026, 24639, 23664, 23173, 22951, 22889, 
    23084, 23639, 24422, 25790, 26533, 21223, 25159, 26585, 26328, 25847, 
    25266, 24745,
  15880, 16071, 21856, 23854, 24989, 24600, 23641, 23106, 22933, 22899, 
    23080, 23535, 24476, 25763, 26635, 21312, 25230, 26566, 26281, 25823, 
    25331, 24854,
  16196, 16396, 22059, 23940, 25041, 24601, 23643, 23135, 22966, 22908, 
    23180, 23518, 24521, 25812, 26771, 21421, 25339, 26587, 26270, 25850, 
    25308, 24741,
  16982, 17195, 22432, 24201, 25096, 24571, 23614, 23183, 22933, 22951, 
    23099, 23573, 24468, 25580, 26660, 21759, 25478, 26618, 26259, 25865, 
    25144, 24676,
  18220, 18407, 23144, 24514, 25151, 24561, 23543, 23114, 22914, 22938, 
    23017, 23589, 24503, 25784, 26541, 22479, 25709, 26597, 26218, 25736, 
    25081, 24409,
  19687, 19786, 24022, 24946, 25208, 24511, 23544, 23113, 22963, 22909, 
    23139, 23665, 24383, 25722, 26991, 23426, 26099, 26626, 26240, 25797, 
    25119, 24531,
  20998, 21028, 24571, 25251, 25274, 24501, 23490, 23117, 22897, 22858, 
    23126, 23706, 24478, 25860, 26934, 24082, 26304, 26572, 26234, 25766, 
    25176, 24646,
  21899, 21915, 24801, 25303, 25325, 24425, 23453, 23087, 22967, 22938, 
    23087, 23712, 24653, 25879, 26907, 24199, 26069, 26558, 26210, 25691, 
    25087, 24514,
  22393, 22455, 24672, 25290, 25229, 24380, 23439, 23064, 22953, 22939, 
    23095, 23664, 24771, 26050, 26881, 23853, 26072, 26436, 26134, 25684, 
    25139, 24588,
  22705, 22820, 24725, 25303, 25234, 24345, 23450, 23108, 22934, 22996, 
    23184, 23739, 24606, 25897, 27081, 23724, 25950, 26515, 26126, 25646, 
    25077, 24514,
  23026, 23151, 25201, 25576, 25290, 24353, 23417, 23097, 22969, 23018, 
    23204, 23667, 24766, 25854, 26922, 24534, 26557, 26562, 26162, 25653, 
    25122, 24702,
  23321, 23429, 25760, 25810, 25361, 24279, 23381, 23064, 22960, 22954, 
    23254, 23646, 24730, 25996, 26902, 25490, 27019, 26610, 26116, 25654, 
    25110, 24522,
  23396, 23499, 25884, 25890, 25333, 24275, 23314, 23034, 22962, 22949, 
    23281, 23739, 24659, 26028, 26800, 25698, 26897, 26493, 26113, 25620, 
    25062, 24429,
  23129, 23259, 25673, 25804, 25224, 24195, 23320, 23047, 22962, 22971, 
    23192, 23757, 24844, 25991, 27279, 25515, 26768, 26481, 26082, 25618, 
    24924, 24325,
  22541, 22654, 25414, 25635, 25158, 24149, 23293, 23042, 22975, 23041, 
    23368, 23841, 24789, 26216, 26921, 24870, 26625, 26423, 26010, 25552, 
    24964, 24302,
  21785, 21753, 25111, 25497, 25066, 24089, 23244, 23007, 22970, 22996, 
    23272, 23867, 24812, 26165, 27457, 23675, 26396, 26435, 25976, 25493, 
    25011, 24412,
  21053, 20825, 25086, 25450, 25020, 24018, 23199, 23039, 22976, 23079, 
    23209, 23942, 24932, 26500, 27116, 23301, 26356, 26285, 25876, 25390, 
    24849, 24268,
  20754, 20414, 25318, 25520, 24940, 23940, 23169, 23023, 22976, 23101, 
    23340, 23847, 25012, 26051, 26674, 23657, 26328, 26225, 25712, 25273, 
    24607, 24109,
  28010, 27958, 27989, 27316, 25889, 24149, 22756, 22266, 22160, 22538, 
    23092, 23675, 24668, 25970, 26661, 28649, 29106, 28135, 27491, 26666, 
    25508, 24461,
  28019, 27981, 28042, 27391, 26042, 24287, 22832, 22284, 22174, 22542, 
    22937, 23668, 24625, 25947, 26793, 28616, 28996, 28031, 27369, 26535, 
    25468, 24415,
  28037, 28037, 27936, 27388, 26070, 24391, 22894, 22316, 22226, 22611, 
    22933, 23679, 24601, 25979, 26943, 28523, 28863, 27875, 27225, 26487, 
    25382, 24282,
  28004, 28054, 27866, 27454, 26189, 24492, 22962, 22408, 22193, 22517, 
    22964, 23579, 24617, 25706, 26726, 28489, 28771, 27779, 27071, 26212, 
    25216, 24107,
  27976, 28056, 27937, 27348, 26271, 24563, 23045, 22441, 22231, 22554, 
    22965, 23537, 24559, 25815, 26580, 28435, 28676, 27697, 26947, 26119, 
    25001, 24026,
  27907, 28010, 27822, 27389, 26318, 24672, 23089, 22479, 22277, 22523, 
    22870, 23584, 24583, 25607, 26979, 28337, 28576, 27642, 26907, 26056, 
    24987, 24073,
  27787, 27888, 27760, 27335, 26339, 24735, 23174, 22521, 22242, 22497, 
    22900, 23567, 24615, 25872, 26663, 28245, 28503, 27335, 26671, 25871, 
    24932, 24032,
  27622, 27709, 27681, 27356, 26374, 24809, 23254, 22575, 22268, 22526, 
    22854, 23522, 24341, 25789, 26883, 28085, 28201, 26959, 26200, 25479, 
    24595, 23965,
  27428, 27505, 27470, 27225, 26319, 24811, 23279, 22580, 22325, 22557, 
    22971, 23487, 24474, 25682, 26804, 27939, 27959, 26760, 26045, 25380, 
    24614, 23959,
  27230, 27309, 27265, 27087, 26291, 24903, 23381, 22656, 22324, 22523, 
    22890, 23496, 24521, 25576, 26691, 27546, 27618, 26447, 25829, 25294, 
    24627, 24080,
  27076, 27150, 26969, 26870, 26212, 24922, 23369, 22676, 22349, 22505, 
    22981, 23584, 24596, 25540, 27029, 27000, 26884, 26157, 25703, 25249, 
    24619, 24092,
  27399, 27347, 26896, 26668, 26010, 24871, 23375, 22601, 22280, 22470, 
    22867, 23474, 24292, 25557, 26663, 26700, 25676, 25577, 25401, 24988, 
    24393, 23817,
  27419, 27332, 26923, 26681, 26028, 24916, 23465, 22622, 22318, 22438, 
    22902, 23400, 24471, 25464, 26513, 26539, 24986, 25159, 25084, 24882, 
    24304, 23864,
  27493, 27381, 26997, 26778, 26122, 24870, 23496, 22672, 22359, 22520, 
    22870, 23440, 24409, 25618, 26726, 26701, 25123, 25202, 25118, 24938, 
    24361, 23917,
  27553, 27442, 27132, 26829, 26196, 24960, 23496, 22698, 22311, 22560, 
    22867, 23410, 24337, 25436, 26554, 26843, 25888, 25519, 25331, 24938, 
    24341, 23970,
  27172, 27204, 26882, 26837, 26323, 25062, 23642, 22824, 22409, 22482, 
    22898, 23432, 24388, 25383, 26751, 26721, 25883, 25578, 25427, 25005, 
    24456, 23873,
  27445, 27360, 27189, 26882, 26284, 25052, 23610, 22792, 22361, 22517, 
    22889, 23419, 24300, 25526, 26498, 26953, 25800, 25476, 25227, 24900, 
    24226, 23809,
  26956, 26992, 26803, 26828, 26338, 25128, 23706, 22867, 22482, 22529, 
    22880, 23471, 24341, 25372, 26482, 26949, 26691, 25981, 25530, 25071, 
    24451, 23742,
  26846, 26877, 26696, 26703, 26341, 25195, 23726, 22904, 22495, 22578, 
    22912, 23545, 24341, 25704, 26562, 26972, 27098, 26306, 25750, 25139, 
    24431, 23895,
  26795, 26822, 26627, 26732, 26323, 25213, 23771, 22960, 22543, 22504, 
    22853, 23487, 24360, 25597, 26388, 26992, 27271, 26422, 25819, 25143, 
    24412, 23795,
  26785, 26830, 26766, 26767, 26361, 25226, 23772, 22982, 22552, 22581, 
    22920, 23366, 24353, 25472, 26606, 27122, 27061, 26292, 25710, 25052, 
    24381, 23795,
  26788, 26867, 26922, 26844, 26330, 25191, 23815, 23029, 22541, 22556, 
    22856, 23495, 24307, 25401, 26794, 27216, 26926, 26197, 25690, 25052, 
    24476, 23728,
  26793, 26903, 26913, 26796, 26382, 25275, 23840, 23072, 22551, 22553, 
    22904, 23412, 24267, 25357, 26749, 27237, 26848, 26212, 25698, 25063, 
    24437, 23746,
  26824, 26932, 26829, 26796, 26379, 25283, 23877, 23065, 22561, 22581, 
    22910, 23433, 24261, 25512, 26500, 27234, 26806, 26179, 25728, 25187, 
    24500, 23779,
  26908, 26964, 26874, 26854, 26401, 25317, 23895, 23076, 22598, 22560, 
    22956, 23396, 24300, 25485, 26758, 27332, 26980, 26256, 25829, 25273, 
    24549, 23857,
  27018, 27028, 27034, 26932, 26466, 25326, 23938, 23108, 22628, 22574, 
    22901, 23455, 24302, 25480, 26419, 27412, 27245, 26490, 25926, 25346, 
    24598, 24021,
  27098, 27115, 26945, 26907, 26419, 25380, 23931, 23098, 22648, 22573, 
    22818, 23388, 24298, 25243, 26577, 27301, 27278, 26484, 26034, 25363, 
    24571, 23900,
  27109, 27188, 26907, 26776, 26385, 25333, 23938, 23087, 22621, 22567, 
    22873, 23486, 24293, 25504, 26613, 27179, 27085, 26432, 25934, 25354, 
    24665, 24033,
  27056, 27185, 26797, 26762, 26318, 25322, 23946, 23152, 22653, 22547, 
    22877, 23401, 24321, 25417, 26261, 27090, 26987, 26369, 25895, 25359, 
    24606, 24006,
  26940, 27081, 26773, 26760, 26281, 25348, 23962, 23152, 22620, 22587, 
    22908, 23437, 24137, 25371, 26478, 27031, 26891, 26337, 25838, 25277, 
    24549, 24026,
  26740, 26868, 26738, 26665, 26284, 25256, 23995, 23143, 22629, 22598, 
    22882, 23311, 24171, 25437, 26503, 27004, 26789, 26340, 25882, 25368, 
    24695, 23887,
  26432, 26556, 26691, 26611, 26255, 25342, 23968, 23151, 22693, 22575, 
    22931, 23386, 24298, 25458, 26361, 26962, 26895, 26344, 25832, 25301, 
    24549, 23994,
  26014, 26145, 26517, 26531, 26205, 25277, 23955, 23155, 22683, 22566, 
    22918, 23360, 24253, 25387, 26169, 26918, 26859, 26253, 25819, 25368, 
    24632, 24001,
  25538, 25665, 26318, 26388, 26160, 25308, 24007, 23179, 22629, 22565, 
    22926, 23389, 24373, 25520, 26481, 26790, 26604, 26246, 25859, 25431, 
    24740, 24074,
  25074, 25207, 26146, 26289, 26109, 25256, 23961, 23205, 22662, 22598, 
    22943, 23343, 24337, 25414, 26143, 26651, 26611, 26134, 25747, 25394, 
    24714, 24101,
  24692, 24862, 25982, 26209, 26023, 25229, 24014, 23179, 22685, 22657, 
    22910, 23294, 24298, 25295, 26390, 26538, 26500, 26076, 25679, 25215, 
    24694, 24041,
  24787, 24867, 26135, 26254, 26016, 25237, 23968, 23121, 22661, 22509, 
    22794, 23283, 24161, 25312, 26525, 26626, 26332, 25904, 25562, 25150, 
    24571, 23984,
  24421, 24624, 25732, 26058, 25968, 25246, 24027, 23220, 22707, 22671, 
    22968, 23359, 24210, 25405, 26369, 26245, 26335, 25893, 25589, 25238, 
    24650, 24136,
  24528, 24651, 25828, 26074, 25999, 25295, 24021, 23253, 22751, 22655, 
    22908, 23353, 24147, 25454, 26425, 26017, 26179, 25881, 25582, 25213, 
    24643, 24051,
  24659, 24690, 25830, 26052, 26029, 25293, 24041, 23242, 22732, 22602, 
    22912, 23315, 24135, 25437, 26899, 25901, 25906, 25869, 25575, 25306, 
    24765, 24106,
  24684, 24667, 25731, 26103, 26040, 25243, 24036, 23273, 22779, 22648, 
    22834, 23387, 24211, 25269, 26263, 26015, 26203, 25932, 25588, 25206, 
    24637, 24020,
  24561, 24533, 25600, 26002, 26004, 25336, 24070, 23244, 22749, 22634, 
    22912, 23304, 24170, 25282, 26810, 25890, 26587, 26069, 25601, 25225, 
    24601, 24102,
  24344, 24325, 25454, 25889, 26003, 25321, 24065, 23316, 22829, 22611, 
    22893, 23340, 24254, 25245, 26325, 25681, 26683, 26101, 25594, 25227, 
    24614, 23970,
  24146, 24134, 25467, 25907, 25965, 25312, 24029, 23258, 22776, 22685, 
    23023, 23368, 24095, 25226, 26624, 25662, 26678, 26113, 25604, 25114, 
    24563, 23976,
  24044, 24041, 25434, 25885, 25961, 25281, 24015, 23230, 22821, 22626, 
    22844, 23339, 24136, 25329, 26241, 25546, 26624, 26113, 25657, 25102, 
    24614, 24015,
  24061, 24061, 25321, 25778, 25971, 25251, 24053, 23250, 22804, 22678, 
    22839, 23358, 24432, 25229, 26569, 25282, 26506, 26132, 25716, 25203, 
    24633, 24076,
  24140, 24146, 25257, 25781, 25931, 25278, 24031, 23249, 22807, 22651, 
    22947, 23346, 24282, 25340, 26715, 25181, 26325, 26059, 25597, 25173, 
    24544, 23933,
  24523, 24398, 25726, 25976, 26019, 25310, 24003, 23236, 22777, 22658, 
    22787, 23346, 24077, 25361, 26420, 25451, 26051, 25781, 25416, 25057, 
    24519, 24017,
  24612, 24500, 25793, 26014, 25988, 25248, 24020, 23182, 22748, 22621, 
    22836, 23316, 24128, 25407, 26029, 25518, 25785, 25485, 25278, 24888, 
    24373, 23930,
  24693, 24604, 25945, 26165, 26082, 25271, 23995, 23191, 22751, 22658, 
    22779, 23336, 24146, 25249, 26445, 25704, 25710, 25312, 25091, 24777, 
    24411, 23943,
  24461, 24538, 25699, 26032, 26037, 25300, 24007, 23268, 22813, 22699, 
    22918, 23394, 24237, 25428, 26421, 25653, 26417, 25921, 25465, 25034, 
    24630, 23929,
  24471, 24577, 25779, 26037, 26068, 25329, 24026, 23273, 22818, 22682, 
    22935, 23422, 24128, 25316, 26381, 25672, 26535, 25953, 25539, 25081, 
    24540, 23976,
  24405, 24537, 25663, 25987, 26024, 25294, 24056, 23291, 22821, 22701, 
    22876, 23292, 24219, 25204, 26644, 25574, 26523, 26106, 25617, 25070, 
    24529, 23978,
  24230, 24381, 25588, 25986, 26032, 25254, 24041, 23307, 22849, 22681, 
    22968, 23361, 24214, 25335, 26606, 25555, 26662, 26209, 25752, 25185, 
    24586, 24044,
  23924, 24104, 25468, 25923, 26006, 25272, 24055, 23292, 22831, 22734, 
    22883, 23386, 24269, 25408, 26563, 25468, 26756, 26346, 25814, 25259, 
    24631, 24072,
  23450, 23674, 25240, 25786, 25937, 25257, 24051, 23304, 22793, 22721, 
    22889, 23320, 24230, 25400, 26407, 25177, 26750, 26524, 25962, 25396, 
    24643, 24098,
  22747, 23009, 25089, 25649, 25865, 25237, 24003, 23282, 22860, 22648, 
    22986, 23336, 24289, 25468, 26415, 24919, 26700, 26688, 26029, 25504, 
    24733, 24172,
  21748, 22022, 24610, 25331, 25744, 25198, 24015, 23264, 22852, 22734, 
    22953, 23396, 24146, 25457, 26539, 24465, 26608, 26801, 26175, 25473, 
    24810, 24093,
  20443, 20739, 23500, 24685, 25479, 25102, 24006, 23271, 22843, 22699, 
    22951, 23398, 24259, 25405, 26710, 23286, 25951, 26770, 26354, 25702, 
    24982, 24227,
  18965, 19298, 22186, 23854, 25135, 25006, 23948, 23289, 22859, 22784, 
    22972, 23436, 24097, 25299, 26707, 21768, 25268, 26717, 26340, 25748, 
    24894, 24314,
  17597, 17961, 21545, 23479, 24975, 25000, 23959, 23255, 22886, 22766, 
    23010, 23387, 24368, 25304, 26559, 21096, 25195, 26700, 26322, 25746, 
    24979, 24154,
  16616, 16986, 21639, 23522, 24979, 24963, 23939, 23225, 22909, 22717, 
    22959, 23467, 24242, 25514, 26876, 21398, 25485, 26704, 26387, 25773, 
    25032, 24370,
  16182, 16533, 21785, 23533, 24952, 24960, 23936, 23274, 22868, 22821, 
    22914, 23426, 24394, 25472, 26854, 21604, 25504, 26681, 26388, 25824, 
    25045, 24474,
  16302, 16613, 21727, 23548, 24969, 24949, 23904, 23293, 22880, 22826, 
    22965, 23442, 24203, 25647, 26713, 21526, 25292, 26737, 26505, 25930, 
    25059, 24442,
  16847, 17132, 21746, 23561, 24968, 24902, 23881, 23269, 22854, 22799, 
    23076, 23447, 24424, 25339, 26721, 21439, 25030, 26672, 26409, 25979, 
    25149, 24376,
  17647, 17918, 22035, 23791, 25009, 24873, 23875, 23226, 22837, 22815, 
    22996, 23408, 24202, 25603, 26713, 21707, 25079, 26700, 26495, 25917, 
    25187, 24470,
  18530, 18788, 22617, 24075, 25115, 24937, 23867, 23210, 22883, 22861, 
    23104, 23467, 24360, 25541, 26667, 22326, 25358, 26649, 26450, 25953, 
    25175, 24482,
  19316, 19572, 23216, 24413, 25217, 24883, 23870, 23285, 22908, 22818, 
    23010, 23436, 24329, 25456, 26682, 22960, 25675, 26760, 26450, 25987, 
    25169, 24472,
  19863, 20146, 23512, 24614, 25276, 24906, 23825, 23219, 22848, 22835, 
    22990, 23520, 24250, 25578, 26935, 23376, 25746, 26697, 26525, 25990, 
    25292, 24474,
  20108, 20447, 23476, 24606, 25330, 24872, 23838, 23193, 22885, 22840, 
    23045, 23447, 24433, 25597, 26573, 23376, 25734, 26744, 26467, 25993, 
    25273, 24689,
  20057, 20471, 23314, 24577, 25234, 24852, 23796, 23187, 22916, 22871, 
    23050, 23504, 24388, 25666, 26676, 23175, 25563, 26704, 26460, 25946, 
    25340, 24589,
  19790, 20247, 23152, 24458, 25261, 24814, 23771, 23197, 22876, 22876, 
    23071, 23538, 24450, 25616, 26831, 22893, 25362, 26695, 26420, 25856, 
    25258, 24607,
  19386, 19831, 23053, 24358, 25197, 24831, 23789, 23192, 22897, 22800, 
    23132, 23487, 24369, 25832, 26784, 22757, 25384, 26643, 26391, 25832, 
    25285, 24636,
  18908, 19296, 22872, 24235, 25170, 24789, 23769, 23190, 22954, 22907, 
    23093, 23492, 24312, 25653, 26595, 22457, 25326, 26604, 26328, 25793, 
    25140, 24649,
  18364, 18718, 22598, 24208, 25157, 24759, 23733, 23189, 22912, 22862, 
    23113, 23456, 24525, 25546, 26551, 22197, 25231, 26565, 26246, 25807, 
    25111, 24604,
  17769, 18109, 22442, 24057, 25087, 24717, 23701, 23171, 22913, 22971, 
    23098, 23526, 24450, 25901, 26708, 21911, 25218, 26585, 26253, 25722, 
    25206, 24539,
  17131, 17475, 22133, 23929, 24999, 24697, 23704, 23213, 22923, 22907, 
    23131, 23522, 24401, 25681, 27166, 21588, 25070, 26497, 26176, 25649, 
    25087, 24578,
  16535, 16848, 21940, 23841, 24974, 24662, 23665, 23137, 22942, 22914, 
    23198, 23593, 24427, 25754, 26801, 21357, 25065, 26601, 26250, 25801, 
    25158, 24526,
  16081, 16355, 21874, 23772, 25032, 24624, 23640, 23231, 22952, 22932, 
    23118, 23504, 24528, 25768, 26835, 21260, 25139, 26570, 26307, 25859, 
    25218, 24768,
  15941, 16164, 21970, 23881, 25009, 24666, 23652, 23191, 22995, 22934, 
    23197, 23631, 24535, 25601, 27002, 21336, 25261, 26659, 26274, 25885, 
    25251, 24655,
  16247, 16475, 22137, 23983, 25073, 24617, 23637, 23196, 22970, 23014, 
    23165, 23623, 24400, 25813, 26901, 21557, 25356, 26615, 26298, 25949, 
    25317, 24710,
  17113, 17345, 22548, 24218, 25082, 24587, 23598, 23139, 22969, 22958, 
    23054, 23638, 24643, 25917, 27250, 21975, 25607, 26559, 26197, 25765, 
    25089, 24544,
  18465, 18667, 23273, 24543, 25177, 24551, 23554, 23157, 22938, 22986, 
    23087, 23620, 24525, 25779, 27167, 22768, 25982, 26532, 26129, 25661, 
    25045, 24392,
  20014, 20138, 24115, 25000, 25262, 24532, 23562, 23148, 22973, 23004, 
    23141, 23712, 24585, 25632, 26925, 23721, 26228, 26538, 26150, 25679, 
    25064, 24433,
  21339, 21408, 24682, 25267, 25323, 24532, 23546, 23102, 22930, 22918, 
    23265, 23588, 24608, 26163, 27112, 24279, 26291, 26528, 26150, 25673, 
    25165, 24548,
  22190, 22249, 24836, 25362, 25329, 24442, 23523, 23118, 22956, 23012, 
    23186, 23698, 24522, 25882, 26699, 24301, 26206, 26492, 26067, 25616, 
    25103, 24456,
  22590, 22687, 24808, 25303, 25314, 24410, 23474, 23116, 22966, 23030, 
    23196, 23638, 24636, 25891, 26881, 24034, 26215, 26377, 25982, 25584, 
    24962, 24423,
  22794, 22926, 24823, 25359, 25288, 24394, 23468, 23089, 23008, 22993, 
    23233, 23728, 24707, 25936, 26999, 23919, 26098, 26362, 25919, 25478, 
    24907, 24303,
  23025, 23150, 25193, 25587, 25349, 24383, 23407, 23090, 22970, 22979, 
    23231, 23757, 24766, 26025, 26894, 24597, 26450, 26373, 25997, 25490, 
    24876, 24390,
  23284, 23388, 25688, 25840, 25380, 24329, 23385, 23102, 23014, 22994, 
    23275, 23836, 24723, 25891, 27231, 25551, 26913, 26472, 25957, 25535, 
    24896, 24431,
  23403, 23510, 25850, 25891, 25304, 24246, 23363, 23124, 22967, 23032, 
    23266, 23794, 24782, 26245, 26928, 25768, 26897, 26420, 25934, 25489, 
    24899, 24318,
  23252, 23398, 25695, 25766, 25235, 24208, 23313, 23090, 23010, 23034, 
    23307, 23826, 24869, 26225, 27281, 25401, 26643, 26407, 25972, 25487, 
    24887, 24227,
  22797, 22937, 25424, 25596, 25175, 24149, 23293, 23056, 22994, 23090, 
    23257, 23835, 24904, 25935, 27034, 24841, 26579, 26436, 25983, 25501, 
    24902, 24358,
  22135, 22143, 25151, 25475, 25060, 24108, 23244, 23075, 23012, 23042, 
    23265, 23989, 24853, 26319, 27265, 23819, 26438, 26412, 25976, 25530, 
    24918, 24381,
  21439, 21265, 25131, 25468, 25006, 23978, 23199, 23067, 23015, 23028, 
    23336, 23936, 24811, 26224, 27077, 23546, 26454, 26276, 25912, 25458, 
    24844, 24264,
  21145, 20867, 25336, 25487, 24940, 23910, 23184, 23077, 22983, 23078, 
    23268, 23892, 24846, 26194, 27310, 23826, 26401, 26101, 25676, 25217, 
    24521, 24038 ;

 CLW =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 
    1, 2, 1, 2, 2, 1, 1, 0, 2, 4, 6, 5, 24, 32, 60, 90, 60, 52, 58, 44, 42, 
    25, 27, 34, 46, 23, 27, 37, 70, 74, 83, 62, 31, 29, 5, 2, 1, 2, 1, 1, 3, 
    2, 1, 2, 1, 1, 4, 5, 10, 15, 0, 0, 0, 9, 13, 3, 1, 2, 6, 9, 14, 14, 2, 0, 
    0, 0, 0, 4, 4, 1, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 5, 5, 
    4, 3, 3, 7, 5, 6, 7, 15, 16, 25, 34, 44, 60, 71, 133, 172, 127, 38, 0, 
    109, 101, 132, 140, 129, 102, 0, 0, 87, 72, 98, 102, 37, 23, 8, 4, 2, 2, 
    2, 1, 2, 0, 1, 0, 0, 1, 1, 2, 4, 19, 8, 0, 0, 0, 2, 13, 6, 6, 11, 17, 24, 
    13, 4, 0, 0, 0, 0, 0, 2, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 5, 7, 11, 
    7, 23, 9, 21, 33, 47, 56, 48, 45, 52, 47, 59, 58, 76, 0, 0, 75, 47, 0, 0, 
    0, 0, 0, 127, 0, 0, 0, 0, 138, 0, 0, 0, 0, 1, 2, 2, 2, 1, 1, 0, 1, 1, 1, 
    0, 1, 1, 3, 23, 17, 0, 0, 0, 0, 8, 12, 14, 18, 19, 19, 17, 9, 0, 0, 0, 0, 
    0, 0, 1, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 2, 21, 18, 19, 
    8, 7, 28, 27, 32, 52, 48, 80, 58, 60, 54, 57, 41, 45, 59, 55, 52, 48, 34, 
    46, 0, 43, 53, 0, 43, 52, 83, 0, 0, 0, 0, 0, 0, 1, 0, 2, 2, 3, 1, 0, 0, 
    0, 0, 0, 2, 2, 4, 16, 16, 16, 0, 0, 0, 0, 10, 16, 21, 17, 14, 8, 7, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 18, 26, 52, 36, 9, 4, 7, 
    10, 3, 4, 11, 19, 24, 29, 56, 52, 45, 50, 84, 98, 85, 72, 72, 0, 56, 52, 
    0, 0, 70, 54, 71, 0, 0, 43, 63, 73, 0, 0, 0, 28, 4, 3, 2, 1, 4, 3, 1, 1, 
    1, 0, 2, 2, 6, 12, 15, 13, 16, 16, 4, 1, 0, 0, 14, 20, 21, 1, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 3, 32, 80, 76, 44, 6, 4, 11, 
    10, 14, 15, 19, 33, 31, 30, 46, 54, 0, 0, 0, 0, 0, 0, 0, 0, 0, 55, 0, 0, 
    23, 70, 0, 0, 76, 0, 0, 0, 28, 0, 0, 8, 4, 3, 3, 2, 4, 2, 1, 0, 2, 2, 4, 
    8, 10, 17, 11, 0, 0, 9, 15, 15, 3, 0, 12, 16, 11, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 29, 85, 63, 16, 12, 5, 3, 
    4, 12, 19, 30, 32, 24, 30, 51, 98, 0, 0, 0, 0, 0, 0, 135, 50, 41, 0, 0, 
    0, 0, 0, 0, 0, 0, 44, 66, 39, 31, 23, 5, 3, 1, 2, 3, 1, 4, 6, 9, 6, 8, 
    12, 13, 10, 10, 2, 0, 0, 0, 1, 17, 16, 2, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 7, 8, 24, 82, 26, 16, 13, 26, 20, 
    20, 21, 30, 50, 41, 31, 53, 63, 64, 92, 99, 87, 107, 0, 0, 73, 70, 78, 
    84, 0, 0, 0, 0, 0, 0, 0, 0, 0, 43, 27, 18, 4, 2, 1, 2, 2, 3, 3, 13, 11, 
    13, 13, 6, 11, 10, 0, 0, 0, 0, 0, 0, 5, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 22, 37, 38, 26, 5, 3, 8, 16, 0, 
    20, 24, 24, 27, 35, 32, 44, 44, 43, 45, 45, 64, 55, 45, 60, 54, 46, 38, 
    58, 59, 0, 0, 0, 0, 0, 0, 0, 0, 27, 22, 0, 0, 0, 3, 3, 2, 7, 6, 6, 2, 11, 
    8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 20, 64, 0, 0, 38, 5, 4, 4, 7, 26, 
    16, 26, 26, 36, 26, 39, 34, 35, 30, 40, 44, 41, 49, 48, 0, 0, 43, 32, 27, 
    46, 72, 0, 0, 33, 0, 0, 0, 29, 23, 0, 1, 0, 1, 4, 8, 5, 8, 6, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 2, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 13, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 63, 37, 46, 0, 0, 44, 3, 2, 5, 36, 59, 
    40, 35, 34, 27, 37, 34, 15, 38, 40, 46, 44, 58, 52, 0, 54, 72, 59, 36, 
    22, 27, 23, 21, 0, 0, 0, 0, 24, 28, 0, 0, 4, 5, 4, 6, 9, 7, 5, 0, 0, 1, 
    1, 0, 0, 0, 0, 3, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 2, 1, 1, 1, 3, 0, 0, 0, 
    0, 0, 3, 6, 11, 6, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 22, 0, 0, 0, 0, 101, 0, 36, 12, 3, 24, 38, 
    48, 42, 32, 33, 11, 28, 30, 38, 63, 40, 41, 67, 50, 61, 0, 44, 41, 54, 
    43, 31, 12, 13, 12, 2, 0, 0, 0, 0, 25, 17, 2, 8, 6, 4, 7, 8, 3, 0, 0, 0, 
    6, 4, 1, 0, 1, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 1, 2, 4, 4, 0, 
    0, 0, 2, 4, 7, 0, 5, 0, 0, 0 ;

 ChanSel =
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1 ;

 ChiSqr =
  0.3410087, 0.3307604, 0.5800743, 0.1674626, 0.1668153, 0.1079943, 
    0.08342511, 0.1909405, 0.2576376, 0.3144295, 0.07539679, 0.2733961, 
    0.5056282, 0.220516, 0.1989998, 0.1353211, 0.1205608, 0.1633477, 
    0.3480781, 0.1325126, 0.2021987, 0.1674835, 0.8640745, 0.2424251, 
    0.2817853, 0.3649582, 0.272792, 0.395526, 0.5551806, 0.5424732, 
    0.2746965, 0.5066894, 0.6362348, 0.4662929, 0.2859842, 0.2147542, 
    0.6672184, 0.3115298, 0.5950376, 0.3544348, 0.5977147, 0.564734, 
    0.4380885, 0.877116, 0.939604, 0.5837358, 0.645557, 0.5047864, 0.6557557, 
    0.6199937, 0.4679467, 0.9475748, 0.400856, 0.4506418, 0.3507315, 
    0.515249, 0.9819729, 0.5634837, 0.3864737, 0.5160101, 0.2938403, 
    0.3144885, 0.6664261, 0.8336596, 0.3343315, 0.2603141, 0.2998693, 
    0.392338, 0.3681831, 0.2408642, 0.3473661, 0.2499139, 0.09093209, 
    0.389369, 0.4413282, 0.4803576, 0.8053818, 0.9583057, 0.3037313, 
    0.262645, 0.181754, 0.2265718, 0.1903346, 0.2682983, 0.08928191, 
    0.8366666, 0.5843719, 0.4525873, 0.1476987, 0.5256856, 0.6216576, 
    0.5725862, 0.2179267, 0.5576022, 0.1932068, 0.4880218,
  0.2487198, 0.2274291, 0.2670563, 0.3356853, 0.05032838, 0.1751546, 
    0.1725441, 0.1441175, 0.211063, 0.3623906, 0.2009079, 0.06762255, 
    0.1464961, 0.1140639, 0.2966029, 0.2464705, 0.1060579, 0.1274645, 
    0.3179381, 0.1034358, 0.2211152, 0.9136658, 0.2705435, 0.4700477, 
    0.2816419, 0.1550951, 0.1767931, 0.9532346, 0.1693208, 0.4667548, 
    0.8605856, 0.8716032, 0.6298108, 0.7719715, 0.6740878, 0.9351029, 
    0.5184001, 0.8647678, 0.3334334, 0.9042587, 2.481207, 1.099246, 
    0.4270862, 0.9525622, 2.994859, 0.9743555, 1.217146, 1.356554, 1.086119, 
    0.9679874, 0.672937, 0.5438589, 0.6725301, 0.7066451, 0.8235267, 
    1.932161, 0.3560041, 0.5925255, 0.7200043, 0.8985796, 0.5264898, 
    0.6029441, 0.5103648, 0.4578457, 0.3430835, 0.3875994, 0.4730046, 
    0.4839646, 0.5023093, 0.5883332, 0.2431807, 0.2065058, 0.3279543, 
    0.3497561, 0.4463853, 0.8680984, 0.9408079, 0.4371923, 0.2543337, 
    0.9077011, 0.2730922, 0.4224937, 0.7175792, 0.1779693, 0.5444967, 
    0.5803025, 0.3278425, 0.1305355, 0.1270331, 0.9965083, 0.5191541, 
    0.2168447, 0.1502331, 0.2189644, 0.1583424, 1.437275,
  0.2624639, 0.209255, 0.2041255, 0.1245288, 0.2445842, 0.2880038, 0.1578767, 
    0.1116685, 0.2267376, 0.36308, 0.4614041, 0.1415786, 0.1135967, 
    0.1388902, 0.227397, 0.1087861, 0.1682538, 0.5143331, 0.2538544, 
    0.4358324, 0.2820921, 0.1875498, 0.4249563, 0.7022278, 0.7600772, 
    0.6036837, 0.7497241, 0.5476046, 0.5111867, 0.4587911, 0.9149452, 
    0.8999217, 0.8175668, 0.3408462, 0.8911608, 0.7132674, 0.4798202, 
    0.8417084, 0.9056906, 0.5086643, 0.3574872, 2.876729, 2.715012, 
    0.8049037, 0.5454962, 0.3318811, 0.3546603, 0.4429584, 2.720055, 
    0.8739386, 0.6141013, 0.8133436, 0.4977386, 4.092341, 0.9960549, 
    0.3365884, 0.3613011, 4.132844, 0.3916101, 0.6033747, 0.2377291, 
    0.6871336, 0.2898677, 0.3854759, 0.4267154, 0.6540501, 0.3844507, 
    0.5100314, 0.5498011, 0.1412097, 0.2209756, 0.1325818, 0.5095547, 
    0.3372023, 0.6590672, 0.8783616, 0.885473, 0.8519764, 0.4241572, 
    0.4431671, 0.4416925, 0.1630915, 0.5723556, 0.3448464, 0.8261992, 
    0.6490891, 0.3045781, 0.1751251, 0.1628084, 0.9429195, 0.2722599, 
    0.3076699, 0.121566, 0.1356849, 0.2865823, 0.2993191,
  0.4289174, 0.3074756, 0.327004, 0.1448061, 0.1239522, 0.1891154, 0.1455189, 
    0.2329021, 0.1449638, 0.2758327, 0.331235, 0.3004084, 0.2948388, 
    0.1541007, 0.05314686, 0.1221706, 0.7069755, 0.7131233, 0.240961, 
    0.3089288, 0.4461661, 0.1911051, 0.3609865, 0.9654834, 0.6679736, 
    0.4514959, 0.765912, 0.6975055, 0.6436234, 0.6967793, 0.6634192, 
    0.7797312, 0.8526489, 0.9193165, 0.3832361, 0.8767279, 0.6860806, 
    0.5781011, 0.8258867, 0.8572273, 2.512301, 1.477677, 0.3014882, 2.875033, 
    0.587013, 0.3680428, 0.73206, 0.75735, 1.100092, 1.016538, 2.077009, 
    0.5562431, 0.7034191, 0.4449839, 0.4858085, 0.2412642, 0.2009655, 
    0.5407128, 0.3619806, 0.7515011, 0.6831266, 0.4401459, 0.3383124, 
    0.7855885, 0.6500106, 0.1502917, 0.1644921, 0.3891912, 0.151869, 
    0.3199321, 0.2498037, 0.9309661, 0.4290444, 0.3160453, 0.9955958, 
    0.7702159, 0.953056, 0.5343935, 0.4393618, 0.8808596, 0.2943498, 
    0.1451782, 0.2695672, 0.4434174, 0.6652893, 1.16585, 0.2056985, 
    0.09583572, 0.09662999, 0.699936, 0.4452049, 0.176788, 0.1618346, 
    0.1265426, 0.2081715, 0.6469927,
  0.5708509, 0.1817875, 0.1355664, 0.165492, 0.1990966, 0.1513804, 
    0.09445122, 0.1239384, 0.2209682, 0.5480772, 0.2235256, 0.1905163, 
    0.1090738, 0.06380407, 0.09635577, 0.3285683, 0.287152, 0.3762916, 
    0.5120324, 0.8065276, 0.8251054, 0.4533577, 0.4736635, 0.6253278, 
    0.4649939, 0.410297, 2.245723, 2.518224, 2.891609, 1.940265, 0.9385162, 
    0.5354626, 0.5000904, 0.7870536, 0.8598505, 0.7734089, 0.9005163, 
    0.6718571, 0.7870947, 0.4783077, 2.269106, 3.515119, 0.3641379, 
    0.5997244, 4.196092, 1.251406, 1.652886, 0.327284, 0.37308, 2.330402, 
    1.323316, 3.513116, 0.5407607, 0.6524888, 0.3056167, 2.680382, 1.46551, 
    0.9540825, 0.5850138, 0.4918625, 0.4373985, 0.322357, 0.3854276, 
    0.3340454, 0.5071886, 0.2364666, 0.2961857, 0.2707906, 0.4267897, 
    0.1712546, 0.3517641, 0.3605876, 0.4571287, 0.8139404, 0.5645651, 
    0.8706505, 0.4648038, 0.260773, 0.3954798, 0.5816071, 0.5864158, 
    0.2841685, 0.574359, 0.9564263, 0.7343218, 0.4179757, 0.2046733, 
    0.8375205, 0.5595151, 0.3125552, 0.2320488, 0.7396886, 0.2677845, 
    0.4516799, 0.2632609, 0.6697785,
  0.3234075, 0.1826984, 0.1364108, 0.1992325, 0.1261351, 0.2888993, 
    0.1010053, 0.1870766, 0.2659398, 0.2081252, 0.1110576, 0.1980008, 
    0.1110308, 0.1035332, 0.7257915, 0.3507305, 0.3445808, 3.589616, 
    0.9043314, 0.7757046, 0.749054, 0.3924482, 0.7340338, 0.7194763, 
    0.3771515, 1.404935, 1.322576, 0.9414355, 2.398568, 2.321282, 0.5065342, 
    0.5269349, 0.4756194, 0.9738931, 0.8800686, 0.5610748, 0.3510796, 
    0.9974131, 0.7533638, 0.7976035, 0.8147787, 3.32464, 0.7246785, 
    0.9813065, 1.503634, 3.274842, 0.3302068, 0.6705939, 1.900696, 0.8027739, 
    0.3381067, 0.5265563, 1.068247, 0.2273645, 0.1742296, 1.502233, 
    0.5940241, 0.7615145, 0.7930545, 0.5413692, 0.4960986, 0.4480969, 
    0.2546907, 0.3533059, 0.2748851, 0.1861418, 0.3463679, 0.3403408, 
    0.5958813, 0.6388312, 0.9904503, 0.8030162, 0.787722, 0.2473987, 
    0.2917701, 0.5573324, 0.72931, 0.2120664, 0.3992558, 0.3410524, 
    0.3898554, 0.5105661, 0.5546927, 0.5501403, 0.3560378, 0.1847725, 
    0.7202161, 0.4337215, 0.7179015, 0.8441041, 0.3983652, 0.2344721, 
    0.2625816, 0.4684231, 0.9757569, 0.5116495,
  0.266003, 0.2268357, 0.1080685, 0.1856613, 0.1995644, 0.1631632, 0.1052112, 
    0.08041472, 0.1599439, 0.1655107, 0.142208, 0.1767619, 0.09813928, 
    0.2736124, 0.4443388, 0.2469674, 0.5251527, 1.591633, 0.7479947, 
    1.452884, 0.821849, 0.6602064, 0.4861808, 0.7199245, 0.6998084, 2.004779, 
    0.4796087, 0.5060464, 0.6653001, 0.399753, 0.4680763, 0.9826325, 
    0.4891014, 0.9250421, 0.9030476, 0.3303654, 0.5319878, 0.4208792, 
    1.696582, 0.4214866, 0.3866094, 0.7020645, 0.4752615, 0.5893473, 
    0.5360413, 0.4427237, 0.705687, 0.7485581, 0.9293699, 2.213039, 1.359392, 
    1.949576, 1.064282, 0.3317119, 2.873829, 0.9447594, 0.3345882, 0.8447512, 
    0.3960887, 0.4531606, 0.5529592, 0.6601287, 0.4501008, 0.3243482, 
    0.4635133, 0.7312295, 0.2687261, 0.3101568, 0.5423341, 0.6226862, 
    0.8238766, 0.9177728, 0.9424626, 0.7273085, 0.3320177, 0.4429994, 
    0.1855165, 0.2712454, 0.6239972, 0.1984728, 0.2318886, 0.7604135, 
    0.6370847, 0.2315596, 0.1559043, 0.6812871, 0.3269231, 0.2309686, 
    0.8578448, 0.6255383, 0.5085959, 0.5338969, 0.2367558, 0.39368, 
    0.6187633, 0.3808962,
  0.1324918, 0.1937323, 0.0700197, 0.1719211, 0.2008985, 0.09764045, 
    0.05042368, 0.101939, 0.198457, 0.1389347, 0.1595318, 0.1021407, 
    0.1245487, 0.3272353, 0.7243764, 0.6750623, 0.4948032, 0.7657669, 
    0.3574999, 1.614533, 2.478608, 0.6024316, 0.8530703, 0.6429183, 1.93185, 
    0.7996904, 0.926413, 0.7145543, 0.2121011, 0.3939292, 0.3261561, 
    0.5217506, 0.6670749, 0.680898, 0.7462967, 3.186574, 0.3863196, 
    0.3989066, 0.9042501, 0.7384522, 1.385917, 4.291928, 0.856208, 0.7756369, 
    0.7212195, 0.9451157, 0.5158188, 0.3200873, 0.3592797, 0.4349352, 
    0.6997862, 0.5613999, 0.6808123, 0.3903232, 0.9481636, 0.9558565, 
    0.3819235, 0.7260937, 0.2382852, 0.2110325, 0.3126152, 0.5656889, 
    0.9945585, 0.3525492, 0.4013632, 0.388853, 0.6891691, 0.4490189, 
    0.7929381, 0.9153424, 0.4674814, 0.9338464, 0.8248432, 0.3539806, 
    0.1052167, 0.1537486, 0.9723231, 0.5385565, 0.7950993, 0.5302549, 
    0.5633033, 0.9951435, 0.6064986, 0.1179393, 0.2613465, 0.2724365, 
    0.264237, 0.2158905, 0.8345357, 0.6564946, 0.2943406, 0.2561976, 
    0.1115318, 0.2160623, 0.5097764, 0.7382724,
  0.1535462, 0.1514977, 0.137351, 0.1190665, 0.1543555, 0.1129074, 
    0.09212694, 0.2840619, 0.1112942, 0.1612339, 0.1406817, 0.9678784, 
    0.3324656, 0.4459544, 0.5260304, 0.883984, 0.3606611, 0.5487729, 
    0.5054317, 0.7751378, 0.8663262, 2.335251, 0.3477467, 3.71834, 0.6329384, 
    0.2837546, 0.2637995, 0.1138478, 0.2467372, 0.3089893, 0.2167469, 
    0.1988744, 0.3115418, 0.2762701, 0.3827906, 0.9091234, 0.9614425, 
    0.6430118, 0.5738366, 0.7278738, 0.3017604, 0.9824137, 1.167756, 
    0.3526183, 0.930303, 0.3547052, 0.4015174, 0.4714632, 0.5986877, 
    0.6998405, 0.4473198, 0.512659, 0.4711796, 0.4782895, 1.234692, 
    0.8792368, 0.4751217, 0.4016696, 0.2616388, 0.6793832, 0.740679, 
    0.5794782, 0.3315835, 0.7933089, 0.7517762, 0.8961377, 0.2980828, 
    0.6671999, 0.6644288, 0.9918033, 0.4471029, 0.8880211, 0.5726717, 
    0.4656965, 0.9188303, 0.8513746, 0.4099633, 0.425854, 0.9439049, 
    0.6029993, 0.3949118, 0.6468663, 0.6155809, 0.1059751, 0.393473, 
    0.279485, 0.8177573, 0.8182267, 0.4716505, 0.210397, 0.2409094, 
    0.1155658, 0.09680921, 0.4125607, 0.3383168, 0.7118473,
  0.4371036, 0.09061962, 0.07627168, 0.1470895, 0.2559217, 0.0622732, 
    0.09139943, 0.1133466, 0.09783449, 0.2654724, 0.621172, 0.4352602, 
    0.1894954, 0.4134946, 0.8183704, 0.3579436, 0.3326386, 0.4316041, 
    0.8141223, 0.1437975, 0.3362018, 0.7328129, 0.3504737, 0.1746008, 
    0.343087, 0.3542572, 0.5436535, 0.2016757, 0.271239, 0.2312961, 
    0.1410555, 0.1129782, 0.2102864, 0.1456408, 0.5865838, 0.6523106, 
    0.6816663, 0.7285075, 0.4339957, 0.5296426, 0.7175869, 0.3037428, 
    0.7787312, 3.640078, 0.3299085, 0.2136239, 1.372227, 0.2741688, 
    0.7551256, 0.4142375, 0.4477501, 0.2872797, 0.2512057, 3.834157, 
    1.308594, 0.448681, 0.5586855, 0.7699007, 0.4438873, 0.9210193, 
    0.7711826, 0.2630808, 0.2888422, 0.2106326, 0.9249786, 1.16522, 
    0.9830437, 0.9495706, 0.6315731, 0.4649216, 0.2354532, 0.360787, 
    0.7733202, 0.5578566, 0.7487851, 0.4326542, 0.4398123, 0.4821829, 
    0.3736224, 0.1421388, 0.3618409, 0.8497465, 0.08521672, 0.06368814, 
    0.4013191, 0.8827225, 0.169713, 0.6967319, 0.409044, 0.2683324, 
    0.1654734, 0.588647, 0.1077542, 0.1954596, 0.3691869, 0.4209514,
  0.1894454, 0.1760956, 0.1285456, 0.08760575, 0.2331225, 0.09320045, 
    0.188126, 0.125982, 0.04302614, 0.154004, 0.3251756, 0.9498312, 
    0.6728074, 0.9523958, 2.643786, 0.8921679, 0.6436291, 0.5998636, 
    0.5695546, 0.4678499, 0.6893415, 0.4030681, 0.7657747, 0.7131853, 
    0.1916575, 0.3463598, 0.3053177, 0.134967, 0.1607937, 0.5687605, 
    0.1722761, 0.1268871, 0.125168, 0.7060817, 0.6271101, 0.3055457, 
    0.5381942, 0.6638797, 2.188019, 0.6463093, 0.6690455, 0.2725076, 
    0.7270026, 0.3020712, 0.8994232, 0.2164283, 0.3977772, 0.4827252, 
    0.3804945, 0.5026218, 0.3418073, 0.1068917, 0.2124953, 2.976359, 
    0.7253647, 0.9031618, 0.3903075, 0.432441, 0.5875769, 0.821734, 
    0.4169648, 0.5505193, 0.4152824, 0.4095642, 0.7120057, 0.224758, 
    0.265657, 0.4962872, 0.1713264, 0.1958164, 0.374347, 0.5768381, 
    0.9688936, 0.3536797, 0.9426571, 0.9983849, 0.3361639, 0.9830844, 
    0.2941018, 0.1889163, 0.3644686, 0.5452048, 0.2721008, 0.1274139, 
    0.4146532, 0.4703127, 0.7312475, 0.4887799, 0.3306941, 0.4709934, 
    0.4324805, 0.1958379, 0.3444948, 0.1443973, 0.3985171, 0.5493177,
  0.3222842, 0.1200974, 0.1162428, 0.1991792, 0.08836729, 0.248246, 
    0.04344666, 0.1136254, 0.6150342, 0.2881329, 0.5272898, 0.2908124, 
    0.6781707, 0.5041931, 0.3075964, 2.724635, 0.2677544, 0.4675604, 
    0.2307717, 0.6475306, 0.218904, 0.127983, 0.2639694, 0.3565804, 
    0.1786332, 0.4314929, 0.7141729, 0.09321578, 0.1144331, 0.2073237, 
    0.3164083, 0.2143066, 0.24299, 0.2609367, 0.3849675, 0.7911157, 
    0.3881373, 0.4100526, 1.006423, 2.822324, 0.83182, 0.9456037, 1.076204, 
    1.591026, 1.114764, 2.671303, 4.67585, 0.2987558, 0.2827561, 0.4961706, 
    0.7650611, 0.9211636, 3.839894, 0.9747463, 0.4015909, 0.8236684, 
    0.4829502, 0.9745503, 0.5416569, 1.768602, 1.174336, 0.6966844, 
    0.6709877, 0.2531933, 0.508689, 0.8160681, 0.4177035, 0.3749397, 
    0.2519612, 0.5416024, 0.8669169, 0.4803922, 0.5929049, 0.4274198, 
    0.5318518, 0.7820568, 0.843772, 0.8488976, 0.4397143, 0.2047727, 
    0.2089693, 0.3590935, 0.3301047, 0.09180469, 0.3234492, 0.4371753, 
    0.6970016, 0.9195036, 0.4721045, 0.2985741, 0.4847079, 0.9856139, 
    0.4702559, 0.2294358, 0.4022827, 0.7356871 ;

 CldBase =
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888 ;

 CldThick =
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888 ;

 CldTop =
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888 ;

 Emis =
  8861, 8964, 9106, 9106, 9106, 9105, 9106, 9106, 9106, 9105, 9105, 9105, 
    9105, 9105, 9105, 9073, 9097, 9097, 9097, 9097, 9097, 9097,
  8840, 8940, 9076, 9079, 9081, 9082, 9085, 9086, 9087, 9090, 9090, 9090, 
    9090, 9090, 9090, 9072, 9210, 9210, 9210, 9210, 9210, 9210,
  8949, 9047, 9134, 9135, 9136, 9137, 9138, 9139, 9139, 9141, 9141, 9141, 
    9141, 9141, 9141, 9127, 9198, 9198, 9197, 9197, 9198, 9198,
  8940, 9035, 9079, 9079, 9079, 9079, 9080, 9080, 9080, 9080, 9080, 9080, 
    9080, 9080, 9080, 9071, 9094, 9094, 9094, 9094, 9094, 9094,
  8959, 9053, 9052, 9054, 9055, 9056, 9058, 9059, 9060, 9062, 9062, 9062, 
    9062, 9062, 9062, 9082, 9146, 9146, 9146, 9146, 9146, 9146,
  8952, 9044, 9038, 9041, 9043, 9044, 9047, 9048, 9049, 9052, 9052, 9052, 
    9052, 9052, 9052, 9070, 9169, 9169, 9169, 9169, 9169, 9169,
  8945, 9045, 8990, 8996, 8999, 9002, 9006, 9008, 9010, 9016, 9016, 9016, 
    9016, 9016, 9016, 9111, 9224, 9224, 9224, 9224, 9224, 9224,
  8875, 8974, 8953, 8958, 8962, 8965, 8969, 8970, 8972, 8978, 8978, 8978, 
    8978, 8978, 8978, 9050, 9187, 9187, 9187, 9187, 9187, 9187,
  8929, 9029, 8979, 8984, 8988, 8990, 8994, 8996, 8998, 9003, 9003, 9003, 
    9003, 9003, 9003, 9092, 9202, 9202, 9202, 9202, 9202, 9202,
  8966, 9065, 9016, 9019, 9021, 9022, 9025, 9026, 9027, 9030, 9030, 9030, 
    9030, 9030, 9030, 9102, 9146, 9146, 9146, 9146, 9146, 9146,
  9004, 9097, 9031, 9039, 9044, 9048, 9054, 9056, 9059, 9068, 9068, 9068, 
    9068, 9068, 9068, 9157, 9375, 9375, 9375, 9375, 9375, 9375,
  9110, 9204, 9081, 9084, 9087, 9089, 9092, 9094, 9095, 9099, 9099, 9099, 
    9099, 9099, 9099, 9199, 9256, 9256, 9256, 9256, 9256, 9256,
  9073, 9166, 9008, 9009, 9009, 9009, 9010, 9011, 9011, 9011, 9011, 9011, 
    9011, 9011, 9011, 9104, 9040, 9040, 9040, 9040, 9040, 9040,
  8982, 9079, 8913, 8917, 8920, 8922, 8925, 8926, 8927, 8932, 8932, 8932, 
    8932, 8932, 8932, 9065, 9084, 9084, 9084, 9084, 9084, 9084,
  9059, 9156, 9008, 9015, 9020, 9024, 9029, 9031, 9034, 9042, 9042, 9042, 
    9042, 9042, 9042, 9187, 9316, 9316, 9316, 9316, 9316, 9316,
  8973, 9068, 8881, 8889, 8894, 8897, 8902, 8904, 8907, 8915, 8915, 8915, 
    8915, 8915, 8915, 9070, 9192, 9192, 9192, 9192, 9192, 9192,
  8994, 9083, 8879, 8887, 8893, 8898, 8903, 8906, 8909, 8919, 8919, 8919, 
    8919, 8919, 8919, 9064, 9244, 9244, 9244, 9244, 9244, 9244,
  8976, 9071, 8747, 8756, 8763, 8767, 8773, 8776, 8779, 8790, 8790, 8790, 
    8790, 8790, 8790, 9023, 9136, 9136, 9136, 9136, 9136, 9136,
  9015, 9115, 8820, 8827, 8831, 8834, 8838, 8840, 8843, 8849, 8849, 8849, 
    8849, 8849, 8849, 9076, 9087, 9087, 9087, 9087, 9087, 9087,
  9001, 9101, 8879, 8883, 8885, 8887, 8890, 8892, 8893, 8897, 8897, 8897, 
    8897, 8897, 8897, 9073, 9052, 9052, 9052, 9052, 9052, 9052,
  9016, 9115, 8928, 8931, 8932, 8934, 8936, 8937, 8938, 8940, 8940, 8940, 
    8940, 8940, 8940, 9083, 9043, 9043, 9043, 9043, 9043, 9043,
  9027, 9129, 8873, 8877, 8880, 8883, 8886, 8887, 8889, 8894, 8894, 8894, 
    8894, 8894, 8894, 9099, 9069, 9068, 9069, 9069, 9068, 9068,
  9157, 9252, 9041, 9042, 9042, 9042, 9043, 9043, 9043, 9044, 9044, 9044, 
    9044, 9044, 9044, 9173, 9067, 9067, 9066, 9066, 9066, 9066,
  9208, 9295, 9032, 9028, 9026, 9024, 9023, 9022, 9021, 9017, 9017, 9017, 
    9017, 9017, 9017, 9118, 8896, 8896, 8896, 8896, 8896, 8896,
  9145, 9237, 8989, 8988, 8987, 8986, 8986, 8986, 8986, 8984, 8984, 8984, 
    8984, 8984, 8984, 9114, 8948, 8948, 8948, 8948, 8948, 8948,
  8962, 9067, 8875, 8877, 8879, 8880, 8883, 8884, 8885, 8888, 8888, 8888, 
    8888, 8888, 8888, 9060, 8996, 8996, 8996, 8996, 8996, 8996,
  8903, 9010, 8767, 8768, 8770, 8770, 8772, 8773, 8773, 8775, 8775, 8775, 
    8775, 8775, 8775, 8975, 8843, 8843, 8843, 8843, 8843, 8843,
  8827, 8941, 8523, 8530, 8535, 8538, 8543, 8545, 8548, 8555, 8555, 8555, 
    8555, 8555, 8555, 8907, 8822, 8822, 8822, 8822, 8822, 8822,
  8850, 8961, 8430, 8435, 8439, 8442, 8446, 8448, 8450, 8456, 8456, 8456, 
    8456, 8456, 8456, 8839, 8666, 8666, 8666, 8666, 8666, 8666,
  8855, 8962, 8537, 8540, 8542, 8544, 8547, 8548, 8549, 8553, 8553, 8553, 
    8553, 8553, 8553, 8858, 8687, 8687, 8687, 8687, 8687, 8687,
  8924, 9031, 8700, 8705, 8708, 8710, 8714, 8715, 8717, 8722, 8722, 8722, 
    8722, 8722, 8722, 8985, 8900, 8900, 8900, 8900, 8900, 8900,
  8980, 9084, 8742, 8746, 8749, 8751, 8755, 8756, 8758, 8762, 8762, 8762, 
    8762, 8762, 8762, 9018, 8928, 8928, 8928, 8928, 8928, 8928,
  9131, 9230, 8839, 8842, 8844, 8845, 8848, 8849, 8850, 8853, 8853, 8853, 
    8853, 8853, 8853, 9109, 8966, 8966, 8966, 8966, 8966, 8966,
  9084, 9179, 8864, 8866, 8867, 8868, 8870, 8870, 8871, 8873, 8873, 8873, 
    8873, 8873, 8873, 9063, 8947, 8947, 8947, 8947, 8947, 8947,
  9137, 9231, 8967, 8967, 8967, 8967, 8967, 8967, 8967, 8967, 8967, 8967, 
    8967, 8967, 8967, 9114, 8962, 8962, 8962, 8962, 8962, 8962,
  9146, 9236, 9003, 9000, 8999, 8997, 8997, 8996, 8995, 8993, 8993, 8993, 
    8993, 8993, 8993, 9096, 8911, 8911, 8911, 8911, 8911, 8911,
  9185, 9273, 9008, 9005, 9004, 9002, 9002, 9000, 9000, 8996, 8996, 8996, 
    8996, 8996, 8996, 9109, 8902, 8902, 8902, 8902, 8902, 8902,
  9306, 9387, 9082, 9076, 9072, 9069, 9067, 9064, 9062, 9056, 9056, 9056, 
    9056, 9056, 9056, 9145, 8845, 8845, 8845, 8845, 8845, 8845,
  9247, 9333, 8884, 8881, 8879, 8877, 8877, 8876, 8874, 8871, 8871, 8871, 
    8871, 8871, 8871, 9065, 8762, 8762, 8762, 8762, 8762, 8762,
  9166, 9257, 8764, 8763, 8762, 8762, 8762, 8762, 8762, 8760, 8760, 8760, 
    8760, 8760, 8760, 9012, 8730, 8730, 8730, 8730, 8730, 8730,
  9125, 9218, 8715, 8715, 8715, 8715, 8716, 8716, 8716, 8715, 8715, 8715, 
    8715, 8715, 8715, 8981, 8715, 8715, 8715, 8715, 8715, 8715,
  9305, 9384, 8877, 8874, 8872, 8870, 8870, 8869, 8868, 8865, 8865, 8865, 
    8865, 8865, 8865, 9062, 8767, 8767, 8767, 8767, 8767, 8767,
  9346, 9421, 8960, 8956, 8954, 8952, 8951, 8950, 8948, 8944, 8944, 8944, 
    8944, 8944, 8944, 9097, 8815, 8815, 8815, 8815, 8815, 8815,
  9329, 9403, 8948, 8943, 8939, 8936, 8934, 8932, 8930, 8924, 8924, 8924, 
    8924, 8924, 8924, 9056, 8725, 8725, 8725, 8725, 8725, 8725,
  9270, 9346, 8931, 8926, 8922, 8919, 8917, 8916, 8914, 8908, 8908, 8908, 
    8908, 8908, 8908, 9026, 8717, 8717, 8717, 8717, 8717, 8717,
  9289, 9363, 9000, 8995, 8991, 8988, 8986, 8985, 8983, 8977, 8977, 8977, 
    8977, 8977, 8977, 9062, 8787, 8787, 8787, 8787, 8787, 8787,
  9491, 9555, 9320, 9307, 9299, 9292, 9287, 9282, 9278, 9264, 9264, 9264, 
    9264, 9264, 9264, 9207, 8814, 8814, 8814, 8814, 8814, 8814,
  9429, 9498, 9176, 9166, 9158, 9153, 9148, 9145, 9141, 9129, 9129, 9129, 
    9129, 9129, 9129, 9148, 8751, 8751, 8751, 8751, 8751, 8751,
  9407, 9474, 9151, 9139, 9132, 9126, 9121, 9117, 9113, 9101, 9101, 9101, 
    9101, 9101, 9101, 9109, 8701, 8701, 8701, 8701, 8701, 8701,
  9301, 9377, 8969, 8964, 8961, 8958, 8956, 8954, 8953, 8947, 8947, 8947, 
    8947, 8947, 8947, 9067, 8765, 8765, 8765, 8765, 8765, 8765,
  9561, 9625, 9253, 9239, 9230, 9222, 9216, 9212, 9207, 9192, 9192, 9192, 
    9192, 9192, 9192, 9200, 8697, 8697, 8697, 8697, 8697, 8697,
  9344, 9419, 9049, 9038, 9031, 9025, 9020, 9017, 9013, 9001, 9001, 9001, 
    9001, 9001, 9001, 9064, 8611, 8611, 8611, 8611, 8611, 8611,
  9227, 9305, 8985, 8978, 8974, 8971, 8968, 8966, 8964, 8957, 8957, 8957, 
    8957, 8957, 8957, 9030, 8736, 8736, 8736, 8736, 8736, 8736,
  9008, 9098, 8764, 8761, 8759, 8758, 8757, 8756, 8755, 8753, 8753, 8753, 
    8753, 8753, 8753, 8901, 8666, 8666, 8666, 8666, 8666, 8666,
  8754, 8859, 8556, 8556, 8556, 8556, 8557, 8557, 8557, 8557, 8557, 8557, 
    8557, 8557, 8557, 8764, 8565, 8565, 8565, 8565, 8565, 8565,
  8543, 8665, 8298, 8301, 8304, 8305, 8308, 8309, 8310, 8314, 8314, 8314, 
    8314, 8314, 8314, 8640, 8447, 8447, 8447, 8447, 8447, 8447,
  8542, 8662, 8175, 8176, 8177, 8178, 8180, 8181, 8181, 8183, 8183, 8183, 
    8183, 8183, 8183, 8552, 8252, 8252, 8252, 8252, 8252, 8252,
  8799, 8906, 8551, 8550, 8549, 8549, 8549, 8549, 8549, 8548, 8548, 8548, 
    8548, 8548, 8548, 8787, 8526, 8526, 8526, 8526, 8526, 8526,
  8847, 8950, 8579, 8578, 8577, 8576, 8577, 8576, 8576, 8574, 8574, 8574, 
    8574, 8574, 8574, 8805, 8536, 8536, 8536, 8536, 8536, 8536,
  8877, 8982, 8841, 8841, 8841, 8841, 8842, 8842, 8842, 8842, 8842, 8842, 
    8842, 8842, 8842, 8973, 8859, 8859, 8859, 8859, 8859, 8859,
  9109, 9219, 9143, 9145, 9147, 9148, 9150, 9151, 9152, 9154, 9154, 9154, 
    9154, 9154, 9154, 9292, 9251, 9251, 9251, 9251, 9251, 9251,
  9308, 9410, 9254, 9257, 9259, 9261, 9263, 9264, 9265, 9268, 9268, 9268, 
    9268, 9268, 9268, 9423, 9382, 9382, 9382, 9382, 9382, 9382,
  9362, 9448, 9225, 9222, 9221, 9219, 9219, 9218, 9217, 9215, 9215, 9215, 
    9215, 9215, 9215, 9301, 9135, 9135, 9135, 9135, 9135, 9135,
  9361, 9444, 9135, 9134, 9134, 9133, 9134, 9133, 9133, 9132, 9132, 9132, 
    9132, 9132, 9132, 9260, 9105, 9105, 9105, 9105, 9105, 9105,
  9442, 9526, 9258, 9257, 9257, 9256, 9257, 9257, 9257, 9256, 9256, 9256, 
    9256, 9256, 9256, 9371, 9242, 9242, 9242, 9242, 9242, 9242,
  9359, 9441, 9188, 9183, 9180, 9177, 9175, 9174, 9172, 9167, 9167, 9167, 
    9167, 9167, 9167, 9239, 8997, 8997, 8997, 8997, 8997, 8997,
  9313, 9398, 9131, 9128, 9125, 9123, 9123, 9121, 9120, 9116, 9116, 9116, 
    9116, 9116, 9116, 9215, 8995, 8995, 8995, 8995, 8995, 8995,
  9305, 9392, 9131, 9132, 9133, 9133, 9134, 9134, 9135, 9136, 9136, 9136, 
    9136, 9136, 9136, 9266, 9172, 9172, 9172, 9172, 9172, 9172,
  9284, 9370, 9071, 9068, 9066, 9064, 9064, 9063, 9062, 9058, 9058, 9058, 
    9058, 9058, 9058, 9177, 8951, 8951, 8951, 8951, 8951, 8951,
  9388, 9475, 9136, 9135, 9134, 9134, 9134, 9134, 9134, 9133, 9133, 9133, 
    9133, 9133, 9133, 9292, 9109, 9108, 9109, 9109, 9108, 9108,
  9361, 9446, 9137, 9139, 9140, 9141, 9143, 9144, 9145, 9147, 9147, 9147, 
    9147, 9147, 9147, 9301, 9230, 9230, 9230, 9230, 9230, 9230,
  9405, 9495, 9230, 9223, 9218, 9215, 9212, 9209, 9207, 9199, 9199, 9199, 
    9199, 9199, 9199, 9297, 8947, 8947, 8947, 8947, 8946, 8947,
  9023, 9132, 9094, 9090, 9087, 9085, 9084, 9083, 9081, 9077, 9077, 9077, 
    9077, 9077, 9077, 9152, 8947, 8947, 8947, 8947, 8947, 8947,
  8452, 8601, 8793, 8801, 8807, 8812, 8817, 8820, 8823, 8833, 8833, 8833, 
    8833, 8833, 8833, 9022, 9164, 9164, 9164, 9164, 9164, 9164,
  7727, 7901, 7811, 7829, 7841, 7851, 7861, 7867, 7873, 7893, 7893, 7893, 
    7893, 7893, 7893, 8364, 8565, 8565, 8565, 8565, 8565, 8565,
  7619, 7820, 7008, 7037, 7057, 7072, 7089, 7099, 7109, 7141, 7141, 7141, 
    7141, 7141, 7141, 8166, 8219, 8219, 8219, 8219, 8219, 8219,
  7588, 7527, 6399, 6440, 6469, 6490, 6511, 6524, 6539, 6583, 6583, 6583, 
    6583, 6583, 6583, 7585, 8083, 8083, 8083, 8083, 8083, 8083,
  7794, 7811, 7072, 7104, 7127, 7144, 7160, 7171, 7183, 7218, 7218, 7218, 
    7218, 7218, 7218, 7946, 8413, 8413, 8413, 8413, 8413, 8413,
  7912, 8074, 7796, 7809, 7819, 7826, 7833, 7838, 7843, 7857, 7857, 7857, 
    7857, 7857, 7857, 8354, 8355, 8355, 8355, 8355, 8355, 8355,
  8248, 8405, 8580, 8590, 8597, 8603, 8609, 8612, 8616, 8627, 8627, 8627, 
    8627, 8627, 8627, 8861, 9013, 9013, 9013, 9013, 9013, 9013,
  8806, 8930, 8950, 8953, 8955, 8957, 8960, 8961, 8962, 8966, 8966, 8966, 
    8966, 8966, 8966, 9113, 9101, 9101, 9101, 9101, 9101, 9101,
  9054, 9161, 9043, 9047, 9050, 9052, 9055, 9057, 9058, 9063, 9063, 9063, 
    9063, 9063, 9063, 9221, 9230, 9230, 9230, 9230, 9230, 9230,
  8942, 9056, 8954, 8957, 8958, 8960, 8962, 8963, 8964, 8967, 8967, 8967, 
    8967, 8967, 8967, 9129, 9070, 9070, 9070, 9070, 9070, 9070,
  8734, 8861, 8919, 8923, 8926, 8928, 8931, 8933, 8934, 8939, 8939, 8939, 
    8939, 8939, 8939, 9084, 9104, 9104, 9104, 9104, 9104, 9104,
  8329, 8485, 8718, 8724, 8728, 8731, 8735, 8736, 8738, 8745, 8745, 8745, 
    8745, 8745, 8745, 8920, 8964, 8964, 8964, 8964, 8964, 8964,
  8045, 8198, 8389, 8396, 8401, 8405, 8409, 8412, 8414, 8422, 8422, 8422, 
    8422, 8422, 8422, 8604, 8693, 8693, 8693, 8693, 8693, 8693,
  7721, 7894, 7834, 7852, 7864, 7874, 7884, 7890, 7897, 7917, 7917, 7917, 
    7917, 7917, 7917, 8371, 8597, 8597, 8597, 8597, 8597, 8597,
  7754, 7925, 7626, 7642, 7652, 7660, 7669, 7675, 7680, 7697, 7697, 7697, 
    7697, 7697, 7697, 8251, 8276, 8276, 8276, 8276, 8276, 8276,
  7370, 7566, 7544, 7557, 7567, 7574, 7580, 7584, 7589, 7604, 7604, 7604, 
    7604, 7604, 7604, 7899, 8092, 8092, 8092, 8092, 8092, 8092,
  7113, 7400, 7603, 7614, 7622, 7627, 7633, 7636, 7640, 7652, 7652, 7652, 
    7652, 7652, 7652, 7963, 8049, 8049, 8049, 8049, 8049, 8049,
  6682, 7037, 7432, 7441, 7448, 7453, 7457, 7460, 7463, 7473, 7473, 7473, 
    7473, 7473, 7473, 7766, 7801, 7801, 7801, 7801, 7801, 7801,
  6194, 6466, 7130, 7160, 7182, 7198, 7214, 7224, 7236, 7270, 7270, 7270, 
    7270, 7270, 7270, 7550, 8328, 8434, 8434, 8434, 8434, 8434,
  5602, 5841, 6544, 6574, 6595, 6611, 6626, 6636, 6648, 6682, 6682, 6682, 
    6682, 6682, 6682, 6911, 7823, 7942, 7942, 7942, 7942, 7942,
  5331, 5573, 6424, 6455, 6477, 6493, 6509, 6519, 6531, 6566, 6566, 6566, 
    6566, 6566, 6566, 6675, 7744, 7865, 7865, 7865, 7865, 7865,
  5534, 5792, 6575, 6607, 6629, 6646, 6662, 6673, 6685, 6721, 6721, 6721, 
    6721, 6721, 6721, 6923, 7897, 8015, 8015, 8015, 8015, 8015,
  5463, 5725, 6096, 6121, 6139, 6152, 6165, 6173, 6182, 6209, 6209, 6209, 
    6209, 6209, 6209, 6396, 7129, 7129, 7129, 7129, 7129, 7129,
  8873, 8978, 9075, 9076, 9076, 9077, 9078, 9078, 9079, 9080, 9080, 9080, 
    9080, 9080, 9080, 9086, 9118, 9118, 9118, 9118, 9118, 9118,
  8838, 8943, 9034, 9037, 9039, 9041, 9043, 9045, 9046, 9049, 9049, 9049, 
    9049, 9049, 9049, 9073, 9178, 9178, 9178, 9178, 9178, 9178,
  8907, 9004, 9136, 9139, 9141, 9142, 9144, 9145, 9146, 9148, 9148, 9148, 
    9148, 9148, 9148, 9112, 9249, 9249, 9249, 9249, 9249, 9249,
  8946, 9044, 9016, 9018, 9018, 9019, 9021, 9021, 9021, 9023, 9023, 9023, 
    9023, 9023, 9023, 9067, 9076, 9076, 9076, 9076, 9076, 9076,
  8915, 9007, 8980, 8983, 8985, 8986, 8988, 8989, 8990, 8993, 8993, 8993, 
    8993, 8993, 8993, 9018, 9100, 9100, 9100, 9100, 9100, 9100,
  9015, 9105, 9083, 9086, 9088, 9089, 9092, 9093, 9094, 9097, 9097, 9097, 
    9097, 9097, 9097, 9120, 9217, 9217, 9217, 9217, 9217, 9217,
  8971, 9065, 9035, 9039, 9042, 9044, 9047, 9048, 9050, 9055, 9055, 9055, 
    9055, 9055, 9055, 9103, 9219, 9219, 9219, 9219, 9219, 9219,
  8983, 9076, 9070, 9077, 9082, 9086, 9090, 9092, 9095, 9103, 9103, 9103, 
    9103, 9103, 9103, 9154, 9367, 9367, 9367, 9367, 9367, 9367,
  8983, 9083, 9018, 9024, 9029, 9032, 9036, 9038, 9041, 9048, 9048, 9048, 
    9048, 9048, 9048, 9154, 9297, 9297, 9297, 9297, 9297, 9297,
  8958, 9055, 8998, 9001, 9004, 9006, 9009, 9010, 9011, 9015, 9015, 9015, 
    9015, 9015, 9015, 9088, 9161, 9161, 9161, 9161, 9161, 9161,
  8975, 9072, 8930, 8936, 8940, 8943, 8946, 8948, 8950, 8957, 8957, 8957, 
    8957, 8957, 8957, 9087, 9177, 9177, 9177, 9177, 9177, 9177,
  9077, 9167, 9023, 9029, 9033, 9036, 9040, 9041, 9043, 9050, 9050, 9050, 
    9050, 9050, 9050, 9152, 9265, 9265, 9265, 9265, 9265, 9265,
  9018, 9111, 8891, 8897, 8901, 8904, 8909, 8910, 8913, 8919, 8919, 8919, 
    8919, 8919, 8919, 9075, 9147, 9147, 9147, 9147, 9147, 9147,
  8987, 9083, 8860, 8868, 8874, 8879, 8884, 8887, 8890, 8899, 8899, 8899, 
    8899, 8899, 8899, 9082, 9223, 9223, 9223, 9223, 9223, 9223,
  9026, 9120, 8946, 8954, 8960, 8964, 8969, 8971, 8974, 8983, 8983, 8983, 
    8983, 8983, 8983, 9128, 9281, 9281, 9281, 9281, 9281, 9281,
  8982, 9075, 8887, 8893, 8898, 8901, 8906, 8908, 8910, 8918, 8918, 8918, 
    8918, 8918, 8918, 9057, 9171, 9171, 9171, 9171, 9171, 9171,
  9059, 9148, 8905, 8911, 8915, 8917, 8921, 8923, 8925, 8932, 8932, 8932, 
    8932, 8932, 8932, 9079, 9150, 9150, 9150, 9150, 9150, 9150,
  9076, 9171, 8862, 8867, 8869, 8872, 8875, 8876, 8878, 8882, 8882, 8882, 
    8882, 8882, 8882, 9082, 9045, 9045, 9045, 9045, 9045, 9045,
  9105, 9209, 8930, 8929, 8928, 8927, 8928, 8928, 8927, 8926, 8926, 8926, 
    8926, 8926, 8926, 9125, 8900, 8900, 8900, 8900, 8900, 8900,
  9029, 9131, 8935, 8938, 8941, 8943, 8945, 8946, 8948, 8952, 8952, 8952, 
    8952, 8952, 8952, 9123, 9094, 9094, 9094, 9094, 9094, 9094,
  9081, 9183, 8992, 8995, 8997, 8999, 9001, 9002, 9003, 9006, 9006, 9006, 
    9006, 9006, 9006, 9169, 9121, 9121, 9121, 9121, 9121, 9121,
  9111, 9206, 9047, 9048, 9048, 9048, 9050, 9050, 9050, 9051, 9051, 9051, 
    9051, 9051, 9051, 9155, 9086, 9086, 9086, 9086, 9086, 9086,
  9227, 9315, 9060, 9056, 9054, 9052, 9051, 9050, 9048, 9044, 9044, 9044, 
    9044, 9044, 9044, 9144, 8917, 8917, 8917, 8917, 8917, 8917,
  9265, 9348, 9038, 9032, 9028, 9025, 9023, 9021, 9019, 9012, 9012, 9012, 
    9012, 9012, 9012, 9103, 8803, 8803, 8803, 8803, 8803, 8803,
  9191, 9279, 9022, 9018, 9016, 9014, 9013, 9012, 9011, 9007, 9007, 9007, 
    9007, 9007, 9007, 9107, 8889, 8889, 8889, 8889, 8889, 8889,
  8971, 9071, 8873, 8872, 8872, 8871, 8872, 8872, 8871, 8870, 8870, 8870, 
    8870, 8870, 8870, 9005, 8847, 8847, 8847, 8847, 8847, 8847,
  8872, 8980, 8740, 8742, 8743, 8744, 8746, 8746, 8747, 8748, 8748, 8748, 
    8748, 8748, 8748, 8947, 8815, 8815, 8815, 8815, 8815, 8815,
  8833, 8940, 8561, 8563, 8564, 8565, 8567, 8567, 8568, 8569, 8569, 8569, 
    8569, 8569, 8569, 8836, 8638, 8638, 8638, 8638, 8638, 8638,
  8949, 9052, 8643, 8643, 8642, 8642, 8642, 8642, 8642, 8641, 8641, 8641, 
    8641, 8641, 8641, 8895, 8628, 8628, 8628, 8628, 8628, 8628,
  8916, 9024, 8680, 8680, 8680, 8680, 8681, 8681, 8681, 8682, 8682, 8682, 
    8682, 8682, 8682, 8927, 8697, 8696, 8697, 8697, 8696, 8696,
  8903, 9009, 8695, 8696, 8696, 8697, 8698, 8698, 8698, 8699, 8699, 8699, 
    8699, 8699, 8699, 8924, 8731, 8731, 8731, 8731, 8731, 8731,
  8985, 9083, 8773, 8771, 8769, 8767, 8767, 8766, 8765, 8762, 8762, 8762, 
    8762, 8762, 8762, 8934, 8677, 8677, 8677, 8677, 8677, 8677,
  9116, 9206, 8760, 8756, 8753, 8751, 8750, 8749, 8748, 8744, 8744, 8744, 
    8744, 8744, 8744, 8948, 8617, 8617, 8617, 8617, 8617, 8617,
  9129, 9220, 8749, 8747, 8746, 8745, 8745, 8744, 8743, 8741, 8741, 8741, 
    8741, 8741, 8741, 8972, 8677, 8677, 8677, 8677, 8677, 8677,
  8946, 9047, 8583, 8583, 8583, 8583, 8584, 8584, 8584, 8583, 8583, 8583, 
    8583, 8583, 8583, 8860, 8585, 8585, 8585, 8585, 8585, 8585,
  9052, 9146, 8798, 8796, 8794, 8793, 8792, 8791, 8790, 8788, 8788, 8788, 
    8788, 8788, 8788, 8965, 8702, 8702, 8702, 8702, 8702, 8702,
  8967, 9068, 8703, 8703, 8704, 8704, 8705, 8705, 8705, 8706, 8706, 8706, 
    8706, 8706, 8706, 8939, 8730, 8730, 8730, 8730, 8730, 8730,
  9149, 9234, 8873, 8867, 8863, 8860, 8858, 8856, 8854, 8847, 8847, 8847, 
    8847, 8847, 8847, 8973, 8639, 8639, 8639, 8639, 8639, 8639,
  8931, 9032, 8630, 8630, 8630, 8630, 8631, 8631, 8631, 8631, 8631, 8631, 
    8631, 8631, 8631, 8877, 8647, 8647, 8647, 8647, 8647, 8647,
  8629, 8745, 8381, 8383, 8385, 8387, 8389, 8390, 8391, 8394, 8394, 8394, 
    8394, 8394, 8394, 8691, 8505, 8505, 8505, 8505, 8505, 8505,
  8497, 8619, 8329, 8332, 8335, 8336, 8339, 8341, 8342, 8346, 8346, 8346, 
    8346, 8346, 8346, 8633, 8484, 8484, 8484, 8484, 8484, 8484,
  8985, 9079, 8662, 8662, 8662, 8662, 8663, 8663, 8663, 8662, 8662, 8662, 
    8662, 8662, 8662, 8885, 8665, 8665, 8665, 8665, 8665, 8665,
  9251, 9330, 8906, 8899, 8894, 8890, 8887, 8885, 8882, 8874, 8874, 8874, 
    8874, 8874, 8874, 9001, 8614, 8614, 8615, 8615, 8614, 8614,
  8792, 8898, 8778, 8781, 8783, 8785, 8787, 8788, 8789, 8792, 8792, 8792, 
    8792, 8792, 8792, 8931, 8906, 8906, 8906, 8906, 8906, 8906,
  8722, 8830, 8418, 8419, 8420, 8420, 8422, 8422, 8423, 8424, 8424, 8424, 
    8424, 8424, 8424, 8703, 8480, 8480, 8480, 8480, 8480, 8480,
  8839, 8939, 8504, 8504, 8504, 8504, 8505, 8505, 8505, 8505, 8505, 8505, 
    8505, 8505, 8505, 8759, 8516, 8516, 8516, 8516, 8516, 8516,
  8435, 8559, 8249, 8252, 8255, 8257, 8259, 8261, 8262, 8266, 8266, 8266, 
    8266, 8266, 8266, 8572, 8411, 8411, 8411, 8411, 8411, 8411,
  8436, 8560, 8254, 8258, 8260, 8262, 8265, 8267, 8268, 8272, 8272, 8272, 
    8272, 8272, 8272, 8575, 8418, 8418, 8418, 8418, 8418, 8418,
  8760, 8865, 8497, 8498, 8499, 8500, 8502, 8502, 8502, 8504, 8504, 8504, 
    8504, 8504, 8504, 8752, 8558, 8558, 8558, 8558, 8558, 8558,
  9008, 9099, 8640, 8639, 8638, 8637, 8638, 8637, 8637, 8635, 8635, 8635, 
    8635, 8635, 8635, 8863, 8597, 8597, 8597, 8597, 8597, 8597,
  8862, 8966, 8830, 8831, 8833, 8834, 8835, 8836, 8837, 8839, 8839, 8839, 
    8839, 8839, 8839, 8967, 8912, 8912, 8912, 8912, 8912, 8912,
  8786, 8895, 8825, 8828, 8830, 8831, 8834, 8835, 8836, 8839, 8839, 8839, 
    8839, 8839, 8839, 8961, 8954, 8954, 8953, 8953, 8954, 8954,
  8787, 8894, 8589, 8590, 8590, 8591, 8592, 8592, 8593, 8593, 8593, 8593, 
    8593, 8593, 8593, 8815, 8630, 8630, 8630, 8630, 8630, 8630,
  8757, 8867, 8550, 8551, 8552, 8553, 8555, 8555, 8556, 8557, 8557, 8557, 
    8557, 8557, 8557, 8801, 8623, 8623, 8623, 8623, 8623, 8623,
  8380, 8508, 8211, 8215, 8218, 8220, 8224, 8225, 8226, 8231, 8231, 8231, 
    8231, 8231, 8231, 8549, 8394, 8394, 8394, 8394, 8394, 8394,
  8266, 8399, 8084, 8089, 8092, 8095, 8099, 8100, 8102, 8107, 8107, 8107, 
    8107, 8107, 8107, 8459, 8298, 8298, 8298, 8298, 8298, 8298,
  8615, 8730, 8278, 8277, 8276, 8275, 8276, 8276, 8275, 8274, 8274, 8274, 
    8274, 8274, 8274, 8589, 8250, 8250, 8250, 8250, 8250, 8250,
  8747, 8860, 8369, 8370, 8371, 8371, 8373, 8373, 8373, 8374, 8374, 8374, 
    8374, 8374, 8374, 8718, 8418, 8418, 8418, 8418, 8418, 8418,
  8863, 8979, 8633, 8632, 8631, 8631, 8632, 8631, 8631, 8630, 8630, 8630, 
    8630, 8630, 8630, 8905, 8613, 8613, 8613, 8613, 8613, 8613,
  8751, 8864, 8652, 8653, 8653, 8653, 8655, 8655, 8655, 8656, 8656, 8656, 
    8656, 8656, 8656, 8855, 8691, 8691, 8691, 8691, 8691, 8691,
  8990, 9099, 8985, 8990, 8994, 8997, 9001, 9003, 9005, 9011, 9011, 9011, 
    9011, 9011, 9011, 9177, 9231, 9231, 9231, 9231, 9231, 9231,
  9177, 9273, 9117, 9117, 9118, 9118, 9120, 9120, 9120, 9121, 9121, 9121, 
    9121, 9121, 9121, 9230, 9156, 9156, 9156, 9156, 9156, 9156,
  9357, 9441, 9233, 9231, 9230, 9228, 9228, 9227, 9227, 9225, 9225, 9225, 
    9225, 9225, 9225, 9298, 9156, 9156, 9156, 9156, 9156, 9156,
  9373, 9457, 9161, 9162, 9162, 9162, 9164, 9164, 9164, 9165, 9165, 9165, 
    9165, 9165, 9165, 9302, 9196, 9196, 9196, 9196, 9196, 9196,
  9424, 9505, 9206, 9203, 9201, 9199, 9198, 9197, 9196, 9192, 9192, 9192, 
    9192, 9192, 9192, 9294, 9080, 9080, 9080, 9080, 9080, 9080,
  9367, 9456, 9166, 9169, 9171, 9172, 9175, 9176, 9177, 9180, 9180, 9180, 
    9180, 9180, 9180, 9348, 9293, 9293, 9293, 9293, 9293, 9293,
  9333, 9421, 9183, 9188, 9191, 9194, 9198, 9199, 9201, 9207, 9207, 9207, 
    9207, 9207, 9207, 9354, 9406, 9406, 9406, 9406, 9406, 9406,
  9242, 9334, 9063, 9068, 9071, 9074, 9077, 9079, 9081, 9086, 9086, 9086, 
    9086, 9086, 9086, 9264, 9278, 9278, 9278, 9278, 9278, 9278,
  9365, 9453, 9158, 9161, 9163, 9164, 9166, 9167, 9168, 9171, 9171, 9171, 
    9171, 9171, 9171, 9334, 9274, 9274, 9274, 9274, 9274, 9274,
  9368, 9455, 9150, 9154, 9157, 9159, 9162, 9163, 9165, 9169, 9169, 9169, 
    9169, 9169, 9169, 9344, 9324, 9324, 9324, 9324, 9324, 9324,
  9334, 9426, 9092, 9093, 9093, 9093, 9094, 9094, 9094, 9095, 9095, 9095, 
    9095, 9095, 9095, 9284, 9119, 9119, 9119, 9119, 9119, 9119,
  9212, 9310, 9116, 9115, 9114, 9113, 9114, 9114, 9113, 9112, 9112, 9112, 
    9112, 9112, 9112, 9241, 9087, 9087, 9087, 9087, 9086, 9087,
  8805, 8934, 8914, 8919, 8922, 8924, 8928, 8930, 8931, 8937, 8937, 8937, 
    8937, 8937, 8937, 9134, 9131, 9131, 9131, 9131, 9131, 9131,
  8137, 8289, 8222, 8236, 8247, 8254, 8263, 8268, 8273, 8290, 8290, 8290, 
    8290, 8290, 8290, 8652, 8849, 8849, 8849, 8849, 8849, 8849,
  7563, 7756, 7305, 7334, 7354, 7370, 7386, 7396, 7406, 7439, 7439, 7439, 
    7439, 7439, 7439, 8245, 8532, 8532, 8532, 8532, 8532, 8532,
  7364, 7575, 6451, 6481, 6503, 6519, 6537, 6548, 6558, 6593, 6593, 6593, 
    6593, 6593, 6593, 7827, 7753, 7753, 7753, 7753, 7753, 7753,
  7179, 7084, 5855, 5903, 5937, 5962, 5988, 6004, 6021, 6074, 6074, 6074, 
    6074, 6074, 6074, 7157, 7858, 7858, 7858, 7858, 7858, 7858,
  7326, 7340, 6504, 6539, 6563, 6582, 6600, 6611, 6624, 6662, 6662, 6662, 
    6662, 6662, 6662, 7513, 7952, 7952, 7952, 7952, 7952, 7952,
  7606, 7792, 7747, 7766, 7779, 7789, 7800, 7807, 7813, 7834, 7834, 7834, 
    7834, 7834, 7834, 8340, 8544, 8544, 8544, 8544, 8544, 8544,
  8094, 8245, 8520, 8527, 8533, 8536, 8541, 8544, 8546, 8555, 8555, 8555, 
    8555, 8555, 8555, 8693, 8839, 8839, 8839, 8839, 8839, 8839,
  8598, 8737, 8920, 8924, 8926, 8929, 8932, 8933, 8934, 8939, 8939, 8939, 
    8939, 8939, 8939, 9067, 9101, 9101, 9101, 9101, 9101, 9101,
  8788, 8916, 8957, 8960, 8963, 8965, 8968, 8969, 8971, 8975, 8975, 8975, 
    8975, 8975, 8975, 9127, 9124, 9124, 9124, 9124, 9124, 9124,
  8639, 8774, 8827, 8832, 8836, 8838, 8842, 8843, 8845, 8850, 8850, 8850, 
    8850, 8850, 8850, 9031, 9040, 9040, 9040, 9040, 9040, 9040,
  8271, 8414, 8536, 8540, 8544, 8546, 8550, 8552, 8553, 8559, 8559, 8559, 
    8559, 8559, 8559, 8728, 8753, 8753, 8753, 8753, 8753, 8753,
  7855, 8015, 8220, 8228, 8233, 8238, 8243, 8245, 8248, 8257, 8257, 8257, 
    8257, 8257, 8257, 8463, 8561, 8561, 8561, 8561, 8561, 8561,
  7683, 7855, 7883, 7893, 7901, 7907, 7913, 7917, 7921, 7933, 7933, 7933, 
    7933, 7933, 7933, 8294, 8348, 8348, 8348, 8348, 8348, 8348,
  7664, 7844, 7419, 7437, 7450, 7460, 7470, 7477, 7483, 7503, 7503, 7503, 
    7503, 7503, 7503, 8176, 8189, 8189, 8189, 8189, 8189, 8189,
  7477, 7626, 7419, 7437, 7450, 7459, 7468, 7474, 7480, 7500, 7500, 7500, 
    7500, 7500, 7500, 7903, 8160, 8160, 8160, 8160, 8160, 8160,
  7207, 7421, 7496, 7509, 7519, 7526, 7533, 7537, 7542, 7557, 7557, 7557, 
    7557, 7557, 7557, 7808, 8056, 8056, 8056, 8056, 8056, 8056,
  7188, 7503, 7749, 7758, 7765, 7770, 7774, 7777, 7780, 7791, 7791, 7791, 
    7791, 7791, 7791, 8129, 8131, 8131, 8131, 8131, 8131, 8131,
  6756, 7105, 7499, 7507, 7513, 7517, 7522, 7524, 7527, 7535, 7535, 7535, 
    7535, 7535, 7535, 7803, 7831, 7831, 7831, 7831, 7831, 7831,
  6336, 6598, 7263, 7292, 7312, 7328, 7342, 7352, 7363, 7395, 7395, 7395, 
    7395, 7395, 7395, 7624, 8391, 8493, 8493, 8493, 8493, 8493,
  5775, 6024, 6681, 6711, 6732, 6748, 6764, 6774, 6785, 6819, 6819, 6819, 
    6819, 6819, 6819, 7102, 7947, 8063, 8063, 8063, 8063, 8063,
  5504, 5762, 6534, 6566, 6588, 6605, 6622, 6632, 6645, 6680, 6680, 6680, 
    6680, 6680, 6680, 6898, 7867, 7987, 7987, 7987, 7987, 7987,
  5670, 5923, 6789, 6820, 6841, 6857, 6873, 6883, 6895, 6928, 6928, 6928, 
    6928, 6928, 6928, 7000, 8029, 8141, 8141, 8141, 8141, 8141,
  5813, 6075, 6988, 7018, 7040, 7056, 7072, 7082, 7093, 7127, 7127, 7127, 
    7127, 7127, 7127, 7150, 8188, 8294, 8294, 8294, 8294, 8294,
  8847, 8953, 9055, 9053, 9052, 9052, 9052, 9051, 9051, 9049, 9049, 9049, 
    9049, 9049, 9049, 9048, 9010, 9010, 9010, 9010, 9010, 9010,
  8864, 8965, 9098, 9100, 9101, 9102, 9103, 9104, 9104, 9106, 9106, 9106, 
    9106, 9106, 9106, 9082, 9172, 9172, 9172, 9172, 9172, 9172,
  8891, 8992, 9101, 9103, 9103, 9104, 9106, 9106, 9107, 9108, 9108, 9108, 
    9108, 9108, 9108, 9098, 9167, 9167, 9167, 9167, 9167, 9167,
  8962, 9057, 9120, 9122, 9123, 9123, 9125, 9125, 9126, 9127, 9127, 9127, 
    9127, 9127, 9127, 9116, 9187, 9187, 9187, 9187, 9187, 9187,
  8981, 9071, 9079, 9081, 9083, 9084, 9087, 9087, 9088, 9091, 9091, 9091, 
    9091, 9091, 9091, 9096, 9197, 9197, 9197, 9197, 9197, 9197,
  9017, 9106, 9079, 9081, 9082, 9084, 9086, 9087, 9087, 9090, 9090, 9090, 
    9090, 9090, 9090, 9110, 9186, 9186, 9186, 9186, 9186, 9186,
  8976, 9065, 9051, 9054, 9056, 9058, 9060, 9062, 9063, 9066, 9066, 9066, 
    9066, 9066, 9066, 9083, 9199, 9199, 9199, 9199, 9199, 9199,
  9000, 9089, 9118, 9123, 9126, 9128, 9131, 9133, 9135, 9140, 9140, 9140, 
    9140, 9140, 9140, 9140, 9318, 9318, 9318, 9318, 9318, 9318,
  8991, 9087, 9026, 9030, 9033, 9036, 9039, 9040, 9042, 9047, 9047, 9047, 
    9047, 9047, 9047, 9120, 9220, 9220, 9220, 9220, 9220, 9220,
  8962, 9058, 8930, 8936, 8940, 8943, 8947, 8948, 8951, 8957, 8957, 8957, 
    8957, 8957, 8957, 9075, 9177, 9177, 9177, 9177, 9177, 9177,
  9008, 9103, 8915, 8919, 8922, 8924, 8927, 8928, 8930, 8934, 8934, 8934, 
    8934, 8934, 8934, 9073, 9094, 9094, 9094, 9094, 9094, 9094,
  9018, 9108, 8953, 8960, 8965, 8968, 8972, 8975, 8977, 8984, 8984, 8984, 
    8984, 8984, 8984, 9095, 9240, 9240, 9240, 9240, 9240, 9240,
  9033, 9126, 8958, 8965, 8969, 8972, 8977, 8979, 8981, 8988, 8988, 8988, 
    8988, 8988, 8988, 9122, 9235, 9235, 9235, 9235, 9235, 9235,
  8990, 9086, 8897, 8906, 8912, 8916, 8922, 8925, 8928, 8937, 8937, 8937, 
    8937, 8937, 8937, 9107, 9266, 9266, 9266, 9266, 9266, 9266,
  9056, 9151, 8957, 8964, 8969, 8972, 8977, 8979, 8982, 8990, 8990, 8990, 
    8990, 8990, 8990, 9150, 9260, 9260, 9260, 9260, 9260, 9260,
  9005, 9100, 8858, 8864, 8868, 8871, 8875, 8877, 8880, 8886, 8886, 8886, 
    8886, 8886, 8886, 9059, 9116, 9116, 9116, 9116, 9116, 9116,
  8990, 9080, 8865, 8869, 8871, 8873, 8876, 8877, 8878, 8882, 8882, 8882, 
    8882, 8882, 8882, 9005, 9024, 9024, 9024, 9024, 9024, 9024,
  9147, 9238, 9123, 9125, 9127, 9128, 9130, 9130, 9131, 9134, 9134, 9134, 
    9134, 9134, 9134, 9209, 9219, 9219, 9219, 9219, 9219, 9219,
  9036, 9140, 8894, 8895, 8895, 8896, 8897, 8897, 8898, 8899, 8899, 8899, 
    8899, 8899, 8899, 9083, 8938, 8938, 8938, 8938, 8938, 8938,
  9011, 9113, 8973, 8974, 8975, 8975, 8977, 8977, 8978, 8979, 8979, 8979, 
    8979, 8979, 8979, 9106, 9030, 9030, 9030, 9030, 9030, 9030,
  9060, 9160, 8992, 8991, 8991, 8991, 8992, 8991, 8991, 8991, 8991, 8991, 
    8991, 8991, 8991, 9114, 8989, 8989, 8989, 8989, 8989, 8989,
  9150, 9239, 9024, 9020, 9017, 9015, 9014, 9013, 9011, 9007, 9007, 9007, 
    9007, 9007, 9007, 9090, 8877, 8877, 8877, 8877, 8877, 8877,
  9238, 9320, 9053, 9047, 9043, 9040, 9038, 9036, 9034, 9027, 9027, 9027, 
    9027, 9027, 9027, 9093, 8820, 8820, 8820, 8820, 8820, 8820,
  9234, 9314, 9042, 9034, 9028, 9024, 9021, 9018, 9015, 9006, 9006, 9006, 
    9006, 9006, 9006, 9053, 8721, 8721, 8721, 8721, 8721, 8721,
  9137, 9222, 8997, 8990, 8985, 8981, 8979, 8976, 8973, 8965, 8965, 8965, 
    8965, 8965, 8965, 9013, 8708, 8708, 8708, 8708, 8708, 8708,
  8931, 9028, 8801, 8797, 8794, 8792, 8791, 8789, 8788, 8783, 8783, 8783, 
    8783, 8783, 8783, 8897, 8644, 8644, 8644, 8644, 8644, 8644,
  8873, 8971, 8537, 8535, 8533, 8532, 8532, 8531, 8531, 8528, 8528, 8528, 
    8528, 8528, 8528, 8761, 8454, 8454, 8454, 8454, 8454, 8454,
  8981, 9077, 8528, 8527, 8526, 8525, 8525, 8525, 8524, 8522, 8522, 8522, 
    8522, 8522, 8522, 8812, 8475, 8475, 8475, 8475, 8475, 8475,
  8812, 8913, 8371, 8369, 8368, 8367, 8367, 8366, 8365, 8363, 8363, 8363, 
    8363, 8363, 8363, 8664, 8300, 8300, 8300, 8300, 8300, 8300,
  8658, 8772, 8397, 8397, 8398, 8399, 8400, 8400, 8401, 8402, 8402, 8402, 
    8402, 8402, 8402, 8685, 8445, 8445, 8445, 8445, 8445, 8445,
  8488, 8612, 8343, 8345, 8347, 8348, 8350, 8351, 8351, 8354, 8354, 8354, 
    8354, 8354, 8354, 8633, 8441, 8441, 8441, 8441, 8441, 8441,
  8553, 8672, 8346, 8346, 8347, 8347, 8348, 8348, 8348, 8349, 8349, 8349, 
    8349, 8349, 8349, 8622, 8374, 8374, 8374, 8374, 8374, 8374,
  8646, 8765, 8376, 8379, 8380, 8382, 8384, 8385, 8385, 8388, 8388, 8388, 
    8388, 8388, 8388, 8710, 8489, 8489, 8489, 8489, 8489, 8489,
  8723, 8835, 8366, 8368, 8369, 8371, 8373, 8374, 8374, 8377, 8377, 8377, 
    8377, 8377, 8377, 8712, 8468, 8468, 8468, 8468, 8468, 8468,
  8838, 8935, 8426, 8424, 8422, 8421, 8421, 8420, 8419, 8416, 8416, 8416, 
    8416, 8416, 8416, 8682, 8335, 8335, 8335, 8335, 8335, 8335,
  8831, 8934, 8387, 8388, 8388, 8389, 8390, 8391, 8391, 8392, 8392, 8392, 
    8392, 8392, 8392, 8722, 8432, 8432, 8432, 8432, 8432, 8432,
  8849, 8950, 8500, 8500, 8499, 8499, 8500, 8500, 8500, 8499, 8499, 8499, 
    8499, 8499, 8499, 8765, 8495, 8495, 8495, 8495, 8495, 8495,
  8930, 9027, 8559, 8558, 8557, 8557, 8557, 8557, 8557, 8555, 8555, 8555, 
    8555, 8555, 8555, 8809, 8531, 8531, 8531, 8531, 8531, 8531,
  8862, 8959, 8572, 8570, 8569, 8568, 8568, 8567, 8566, 8564, 8564, 8564, 
    8564, 8564, 8564, 8769, 8497, 8497, 8497, 8497, 8497, 8497,
  8611, 8729, 8695, 8699, 8701, 8703, 8706, 8707, 8709, 8712, 8712, 8712, 
    8712, 8712, 8712, 8854, 8855, 8855, 8855, 8855, 8855, 8855,
  8592, 8710, 8636, 8639, 8642, 8643, 8646, 8647, 8649, 8652, 8652, 8652, 
    8652, 8652, 8652, 8815, 8792, 8792, 8792, 8792, 8792, 8792,
  8959, 9053, 8694, 8692, 8691, 8690, 8690, 8690, 8689, 8687, 8687, 8687, 
    8687, 8687, 8687, 8873, 8638, 8638, 8638, 8638, 8638, 8638,
  8943, 9036, 8696, 8690, 8685, 8682, 8679, 8677, 8675, 8667, 8667, 8667, 
    8667, 8667, 8667, 8807, 8435, 8435, 8435, 8435, 8435, 8435,
  8549, 8669, 8536, 8540, 8543, 8546, 8549, 8551, 8552, 8557, 8557, 8557, 
    8557, 8557, 8557, 8763, 8739, 8739, 8739, 8739, 8739, 8739,
  8486, 8609, 8513, 8518, 8521, 8524, 8527, 8529, 8531, 8536, 8536, 8536, 
    8536, 8536, 8536, 8738, 8732, 8732, 8732, 8732, 8732, 8732,
  8501, 8624, 8555, 8560, 8563, 8565, 8568, 8569, 8571, 8576, 8576, 8576, 
    8576, 8576, 8576, 8759, 8745, 8745, 8745, 8745, 8745, 8745,
  8507, 8631, 8590, 8594, 8597, 8599, 8602, 8603, 8605, 8609, 8609, 8609, 
    8609, 8609, 8609, 8778, 8772, 8772, 8772, 8772, 8772, 8772,
  8571, 8691, 8674, 8678, 8681, 8683, 8686, 8687, 8689, 8693, 8693, 8693, 
    8693, 8693, 8693, 8835, 8846, 8846, 8846, 8846, 8846, 8846,
  8448, 8571, 8294, 8297, 8299, 8301, 8304, 8305, 8306, 8309, 8309, 8309, 
    8309, 8309, 8309, 8590, 8437, 8437, 8437, 8437, 8437, 8437,
  8684, 8797, 8721, 8724, 8726, 8728, 8730, 8731, 8732, 8736, 8736, 8736, 
    8736, 8736, 8736, 8880, 8858, 8858, 8858, 8858, 8858, 8858,
  8680, 8797, 8747, 8750, 8753, 8755, 8757, 8758, 8760, 8763, 8763, 8763, 
    8763, 8763, 8763, 8911, 8900, 8900, 8900, 8900, 8900, 8900,
  8618, 8739, 8726, 8730, 8733, 8735, 8738, 8739, 8741, 8745, 8745, 8745, 
    8745, 8745, 8745, 8892, 8902, 8902, 8902, 8902, 8902, 8902,
  8526, 8652, 8632, 8637, 8641, 8643, 8647, 8648, 8650, 8656, 8656, 8656, 
    8656, 8656, 8656, 8832, 8852, 8852, 8852, 8852, 8852, 8852,
  8127, 8273, 7937, 7943, 7947, 7950, 7954, 7956, 7958, 7964, 7964, 7964, 
    7964, 7964, 7964, 8382, 8189, 8189, 8189, 8189, 8189, 8189,
  8411, 8543, 8466, 8472, 8477, 8480, 8485, 8487, 8489, 8496, 8496, 8496, 
    8496, 8496, 8496, 8736, 8750, 8750, 8750, 8750, 8750, 8750,
  8315, 8451, 8335, 8342, 8347, 8350, 8355, 8357, 8359, 8367, 8367, 8367, 
    8367, 8367, 8367, 8639, 8630, 8630, 8630, 8630, 8630, 8630,
  8359, 8489, 8324, 8328, 8332, 8334, 8337, 8339, 8341, 8346, 8346, 8346, 
    8346, 8346, 8346, 8606, 8528, 8528, 8528, 8528, 8528, 8528,
  8633, 8767, 8328, 8331, 8333, 8335, 8337, 8338, 8339, 8342, 8342, 8342, 
    8342, 8342, 8342, 8762, 8458, 8458, 8458, 8458, 8458, 8458,
  8715, 8841, 8458, 8461, 8463, 8465, 8467, 8468, 8469, 8473, 8473, 8473, 
    8473, 8473, 8473, 8835, 8598, 8598, 8598, 8598, 8598, 8598,
  8724, 8841, 8567, 8570, 8573, 8574, 8577, 8578, 8579, 8583, 8583, 8583, 
    8583, 8583, 8583, 8846, 8718, 8718, 8718, 8718, 8718, 8718,
  8896, 9007, 8927, 8930, 8933, 8935, 8938, 8940, 8941, 8945, 8945, 8945, 
    8945, 8945, 8945, 9093, 9103, 9103, 9103, 9103, 9103, 9103,
  9123, 9222, 9103, 9104, 9106, 9107, 9108, 9109, 9110, 9112, 9112, 9112, 
    9112, 9112, 9112, 9217, 9186, 9186, 9186, 9186, 9186, 9186,
  9334, 9424, 9192, 9192, 9193, 9193, 9194, 9194, 9194, 9195, 9195, 9195, 
    9195, 9195, 9195, 9321, 9226, 9226, 9226, 9226, 9226, 9226,
  9423, 9506, 9195, 9197, 9199, 9200, 9202, 9202, 9203, 9205, 9205, 9205, 
    9205, 9205, 9205, 9353, 9287, 9287, 9287, 9287, 9287, 9287,
  9498, 9582, 9223, 9228, 9231, 9233, 9236, 9238, 9239, 9244, 9244, 9244, 
    9244, 9244, 9244, 9441, 9418, 9418, 9418, 9418, 9418, 9418,
  9434, 9517, 9210, 9213, 9214, 9215, 9218, 9218, 9219, 9222, 9222, 9222, 
    9222, 9222, 9222, 9371, 9317, 9317, 9317, 9317, 9317, 9317,
  9334, 9419, 9119, 9121, 9123, 9124, 9127, 9127, 9128, 9131, 9131, 9131, 
    9131, 9131, 9131, 9284, 9232, 9232, 9232, 9232, 9232, 9232,
  9333, 9419, 9147, 9152, 9155, 9157, 9161, 9162, 9164, 9169, 9169, 9169, 
    9169, 9169, 9169, 9324, 9351, 9351, 9351, 9351, 9351, 9351,
  9264, 9358, 9039, 9045, 9049, 9052, 9056, 9058, 9060, 9067, 9067, 9067, 
    9067, 9067, 9067, 9287, 9297, 9297, 9297, 9297, 9297, 9297,
  9206, 9303, 9062, 9065, 9068, 9070, 9073, 9074, 9075, 9079, 9079, 9079, 
    9079, 9079, 9079, 9255, 9227, 9227, 9227, 9227, 9227, 9227,
  9086, 9193, 8980, 8980, 8981, 8981, 8983, 8983, 8983, 8984, 8984, 8984, 
    8984, 8984, 8984, 9173, 9025, 9025, 9025, 9025, 9025, 9025,
  8852, 8975, 8946, 8949, 8952, 8953, 8956, 8957, 8959, 8963, 8963, 8963, 
    8963, 8963, 8963, 9129, 9103, 9103, 9103, 9103, 9103, 9103,
  8455, 8607, 8680, 8687, 8691, 8694, 8699, 8701, 8703, 8710, 8710, 8710, 
    8710, 8710, 8710, 8958, 8955, 8955, 8955, 8955, 8955, 8955,
  7984, 8146, 7844, 7860, 7871, 7880, 7890, 7895, 7901, 7919, 7919, 7919, 
    7919, 7919, 7919, 8453, 8535, 8535, 8535, 8535, 8535, 8535,
  7396, 7545, 6960, 6977, 6989, 6999, 7008, 7013, 7021, 7041, 7041, 7041, 
    7041, 7041, 7041, 8218, 7904, 8017, 8017, 8017, 8017, 8017,
  7084, 7058, 5966, 6013, 6046, 6070, 6094, 6110, 6126, 6178, 6178, 6178, 
    6178, 6178, 6178, 7316, 7905, 7905, 7905, 7905, 7905, 7905,
  6958, 6895, 5813, 5865, 5901, 5928, 5954, 5972, 5990, 6046, 6046, 6046, 
    6046, 6046, 6046, 7099, 7945, 7945, 7945, 7945, 7945, 7945,
  7297, 7371, 6838, 6874, 6899, 6917, 6936, 6947, 6960, 6999, 6999, 6999, 
    6999, 6999, 6999, 7712, 8307, 8307, 8307, 8307, 8307, 8307,
  7347, 7537, 7651, 7665, 7674, 7682, 7690, 7695, 7700, 7715, 7715, 7715, 
    7715, 7715, 7715, 8120, 8244, 8244, 8244, 8244, 8244, 8244,
  7716, 7895, 8410, 8426, 8437, 8446, 8455, 8461, 8466, 8484, 8484, 8484, 
    8484, 8484, 8484, 8659, 9097, 9097, 9097, 9097, 9097, 9097,
  8168, 8320, 8564, 8569, 8573, 8575, 8579, 8581, 8583, 8588, 8588, 8588, 
    8588, 8588, 8588, 8730, 8790, 8790, 8790, 8790, 8790, 8790,
  8242, 8385, 8376, 8385, 8392, 8397, 8403, 8406, 8410, 8420, 8420, 8420, 
    8420, 8420, 8420, 8687, 8786, 8786, 8786, 8786, 8786, 8786,
  8054, 8209, 8102, 8115, 8124, 8131, 8139, 8143, 8148, 8162, 8162, 8162, 
    8162, 8162, 8162, 8546, 8656, 8656, 8656, 8656, 8656, 8656,
  7680, 7855, 7778, 7793, 7803, 7811, 7820, 7825, 7830, 7846, 7846, 7846, 
    7846, 7846, 7846, 8300, 8403, 8403, 8403, 8403, 8403, 8403,
  7518, 7700, 7670, 7685, 7695, 7703, 7713, 7718, 7723, 7740, 7740, 7740, 
    7740, 7740, 7740, 8199, 8321, 8321, 8321, 8321, 8321, 8321,
  7482, 7668, 7317, 7335, 7348, 7358, 7369, 7376, 7382, 7403, 7403, 7403, 
    7403, 7403, 7403, 8062, 8113, 8113, 8113, 8113, 8113, 8113,
  7485, 7597, 7222, 7250, 7271, 7286, 7300, 7310, 7320, 7352, 7352, 7352, 
    7352, 7352, 7352, 7942, 8412, 8411, 8411, 8412, 8412, 8411,
  7256, 7376, 7149, 7173, 7190, 7203, 7215, 7223, 7232, 7259, 7259, 7259, 
    7259, 7259, 7259, 7654, 8154, 8154, 8154, 8154, 8154, 8154,
  7138, 7373, 7469, 7483, 7493, 7500, 7507, 7511, 7516, 7531, 7531, 7531, 
    7531, 7531, 7531, 7825, 8037, 8037, 8037, 8037, 8037, 8037,
  7223, 7553, 7835, 7841, 7845, 7848, 7851, 7853, 7855, 7861, 7861, 7861, 
    7861, 7861, 7861, 8171, 8078, 8078, 8078, 8078, 8078, 8078,
  6888, 7253, 7727, 7729, 7730, 7731, 7732, 7732, 7732, 7734, 7734, 7734, 
    7734, 7734, 7734, 7892, 7789, 7789, 7789, 7789, 7790, 7790,
  6423, 6863, 7506, 7511, 7515, 7518, 7521, 7522, 7524, 7530, 7530, 7530, 
    7530, 7530, 7530, 7779, 7721, 7721, 7721, 7721, 7721, 7721,
  5952, 6197, 6943, 6971, 6992, 7007, 7022, 7031, 7043, 7075, 7075, 7075, 
    7075, 7075, 7075, 7222, 8119, 8227, 8227, 8227, 8227, 8227,
  5731, 5968, 6766, 6795, 6815, 6831, 6846, 6855, 6867, 6899, 6899, 6899, 
    6899, 6899, 6899, 6997, 7973, 8085, 8085, 8085, 8085, 8085,
  5703, 5922, 6707, 6734, 6753, 6768, 6782, 6791, 6801, 6832, 6832, 6832, 
    6832, 6832, 6832, 6898, 7880, 7992, 7992, 7992, 7992, 7992,
  5764, 6008, 7049, 7078, 7098, 7113, 7128, 7137, 7148, 7180, 7180, 7180, 
    7180, 7180, 7180, 7018, 8180, 8282, 8282, 8282, 8282, 8282,
  8831, 8937, 9049, 9047, 9045, 9044, 9044, 9043, 9042, 9040, 9040, 9040, 
    9040, 9040, 9040, 9026, 8967, 8967, 8967, 8967, 8967, 8967,
  8810, 8916, 8985, 8984, 8983, 8982, 8982, 8982, 8981, 8980, 8980, 8980, 
    8980, 8980, 8980, 8992, 8938, 8938, 8937, 8937, 8938, 8938,
  8881, 8989, 9027, 9028, 9028, 9028, 9029, 9029, 9029, 9030, 9030, 9030, 
    9030, 9030, 9030, 9082, 9054, 9054, 9054, 9054, 9054, 9054,
  8892, 8990, 9049, 9049, 9049, 9049, 9050, 9050, 9050, 9050, 9050, 9050, 
    9050, 9050, 9050, 9048, 9064, 9064, 9064, 9064, 9064, 9064,
  8936, 9033, 9015, 9016, 9017, 9018, 9020, 9020, 9021, 9022, 9022, 9022, 
    9022, 9022, 9022, 9061, 9084, 9084, 9084, 9084, 9084, 9084,
  9053, 9142, 9156, 9159, 9161, 9163, 9165, 9166, 9167, 9171, 9171, 9171, 
    9171, 9171, 9171, 9172, 9296, 9296, 9296, 9296, 9296, 9296,
  8971, 9065, 8988, 8992, 8995, 8997, 9000, 9001, 9003, 9007, 9007, 9007, 
    9007, 9007, 9007, 9079, 9161, 9161, 9161, 9161, 9161, 9161,
  9031, 9125, 9107, 9111, 9114, 9117, 9120, 9121, 9123, 9128, 9128, 9128, 
    9128, 9128, 9128, 9178, 9308, 9308, 9308, 9308, 9308, 9308,
  8990, 9082, 9029, 9036, 9041, 9045, 9049, 9051, 9054, 9062, 9062, 9062, 
    9062, 9062, 9062, 9131, 9327, 9327, 9327, 9327, 9327, 9327,
  8957, 9053, 8919, 8925, 8929, 8932, 8936, 8938, 8940, 8947, 8947, 8947, 
    8947, 8947, 8947, 9069, 9172, 9172, 9172, 9172, 9172, 9172,
  8980, 9078, 8933, 8938, 8942, 8945, 8949, 8951, 8953, 8959, 8959, 8959, 
    8959, 8959, 8959, 9092, 9171, 9171, 9171, 9171, 9171, 9171,
  8914, 9012, 8865, 8872, 8877, 8880, 8885, 8887, 8890, 8898, 8898, 8898, 
    8898, 8898, 8898, 9040, 9168, 9168, 9168, 9168, 9168, 9168,
  9000, 9101, 8877, 8883, 8887, 8891, 8895, 8897, 8899, 8906, 8906, 8906, 
    8906, 8906, 8906, 9101, 9145, 9145, 9145, 9145, 9145, 9145,
  9030, 9125, 8959, 8967, 8972, 8976, 8981, 8984, 8987, 8995, 8995, 8995, 
    8995, 8995, 8995, 9146, 9292, 9292, 9292, 9292, 9292, 9292,
  9019, 9118, 8950, 8954, 8956, 8958, 8961, 8962, 8963, 8967, 8967, 8967, 
    8967, 8967, 8967, 9107, 9104, 9104, 9104, 9104, 9104, 9104,
  8997, 9101, 8866, 8866, 8867, 8867, 8868, 8868, 8868, 8868, 8868, 8868, 
    8868, 8868, 8868, 9044, 8885, 8885, 8885, 8885, 8885, 8885,
  9092, 9188, 9049, 9048, 9048, 9047, 9048, 9048, 9048, 9047, 9047, 9047, 
    9047, 9047, 9047, 9137, 9031, 9031, 9031, 9031, 9031, 9031,
  9080, 9176, 9049, 9047, 9047, 9046, 9046, 9046, 9045, 9044, 9044, 9044, 
    9044, 9044, 9044, 9126, 9011, 9011, 9011, 9011, 9011, 9011,
  9090, 9192, 8997, 8997, 8997, 8997, 8998, 8998, 8998, 8998, 8998, 8998, 
    8998, 8998, 8998, 9144, 9010, 9010, 9010, 9010, 9010, 9010,
  9040, 9139, 8957, 8956, 8955, 8954, 8955, 8954, 8954, 8953, 8953, 8953, 
    8953, 8953, 8953, 9075, 8923, 8923, 8923, 8923, 8922, 8923,
  9079, 9174, 8973, 8975, 8976, 8977, 8978, 8979, 8980, 8981, 8981, 8981, 
    8981, 8981, 8981, 9113, 9049, 9049, 9049, 9049, 9049, 9049,
  9130, 9217, 8845, 8841, 8839, 8837, 8836, 8835, 8833, 8829, 8829, 8829, 
    8829, 8829, 8829, 8982, 8703, 8703, 8703, 8703, 8703, 8703,
  9219, 9299, 8946, 8940, 8935, 8932, 8930, 8927, 8925, 8918, 8918, 8918, 
    8918, 8918, 8918, 9018, 8690, 8690, 8690, 8690, 8690, 8690,
  9172, 9254, 9011, 9002, 8996, 8991, 8987, 8984, 8981, 8971, 8971, 8971, 
    8971, 8971, 8971, 9006, 8646, 8646, 8646, 8646, 8646, 8646,
  9032, 9125, 8886, 8882, 8879, 8877, 8876, 8874, 8873, 8868, 8868, 8868, 
    8868, 8868, 8868, 8973, 8726, 8726, 8726, 8726, 8726, 8726,
  9015, 9114, 8797, 8797, 8796, 8796, 8796, 8796, 8796, 8795, 8795, 8795, 
    8795, 8795, 8795, 8982, 8775, 8775, 8775, 8775, 8775, 8775,
  8955, 9047, 8522, 8520, 8518, 8517, 8517, 8516, 8515, 8512, 8512, 8512, 
    8512, 8512, 8512, 8772, 8438, 8438, 8438, 8438, 8438, 8438,
  8933, 9027, 8416, 8415, 8413, 8413, 8413, 8412, 8411, 8409, 8409, 8409, 
    8409, 8409, 8409, 8720, 8355, 8355, 8355, 8355, 8355, 8355,
  8861, 8962, 8393, 8393, 8392, 8392, 8393, 8392, 8392, 8391, 8391, 8391, 
    8391, 8391, 8391, 8717, 8377, 8377, 8377, 8377, 8377, 8377,
  8600, 8717, 8311, 8313, 8313, 8314, 8316, 8316, 8317, 8318, 8318, 8318, 
    8318, 8318, 8318, 8633, 8376, 8376, 8376, 8376, 8376, 8376,
  8475, 8607, 8333, 8337, 8340, 8342, 8345, 8347, 8348, 8353, 8353, 8353, 
    8353, 8353, 8353, 8681, 8518, 8518, 8518, 8518, 8518, 8518,
  8146, 8296, 8041, 8048, 8053, 8057, 8061, 8064, 8066, 8074, 8074, 8074, 
    8074, 8074, 8074, 8479, 8349, 8349, 8349, 8349, 8349, 8349,
  8549, 8673, 8168, 8172, 8175, 8177, 8180, 8181, 8183, 8187, 8187, 8187, 
    8187, 8187, 8187, 8603, 8348, 8348, 8348, 8348, 8348, 8348,
  8730, 8842, 8395, 8397, 8399, 8401, 8403, 8404, 8405, 8408, 8408, 8408, 
    8408, 8408, 8408, 8737, 8520, 8520, 8520, 8520, 8520, 8520,
  8737, 8847, 8330, 8332, 8334, 8335, 8338, 8339, 8339, 8342, 8342, 8342, 
    8342, 8342, 8342, 8695, 8444, 8444, 8444, 8444, 8444, 8444,
  8869, 8970, 8444, 8445, 8445, 8446, 8447, 8448, 8448, 8449, 8449, 8449, 
    8449, 8449, 8449, 8764, 8490, 8490, 8490, 8490, 8490, 8490,
  8972, 9069, 8562, 8562, 8562, 8562, 8563, 8563, 8563, 8563, 8563, 8563, 
    8563, 8563, 8563, 8849, 8573, 8573, 8573, 8573, 8573, 8573,
  9112, 9201, 8769, 8767, 8766, 8765, 8765, 8765, 8764, 8762, 8762, 8762, 
    8762, 8762, 8762, 8965, 8712, 8712, 8712, 8712, 8712, 8712,
  8997, 9092, 8666, 8666, 8665, 8665, 8666, 8665, 8665, 8664, 8664, 8664, 
    8664, 8664, 8664, 8894, 8653, 8653, 8653, 8653, 8653, 8653,
  8891, 8986, 8616, 8613, 8610, 8608, 8607, 8605, 8604, 8600, 8600, 8600, 
    8600, 8600, 8600, 8778, 8464, 8464, 8464, 8464, 8464, 8464,
  8813, 8912, 8555, 8551, 8548, 8546, 8546, 8544, 8543, 8539, 8539, 8539, 
    8539, 8539, 8539, 8729, 8412, 8412, 8412, 8412, 8412, 8412,
  8812, 8914, 8590, 8587, 8584, 8583, 8582, 8581, 8579, 8576, 8576, 8576, 
    8576, 8576, 8576, 8760, 8459, 8459, 8459, 8459, 8459, 8459,
  8663, 8773, 8397, 8393, 8391, 8389, 8388, 8387, 8385, 8381, 8381, 8381, 
    8381, 8381, 8381, 8620, 8255, 8255, 8255, 8255, 8255, 8255,
  8707, 8813, 8485, 8481, 8477, 8475, 8474, 8472, 8471, 8465, 8465, 8465, 
    8465, 8465, 8465, 8657, 8308, 8308, 8308, 8308, 8308, 8308,
  8460, 8585, 8468, 8474, 8477, 8480, 8484, 8486, 8488, 8494, 8494, 8494, 
    8494, 8494, 8494, 8713, 8710, 8710, 8710, 8710, 8710, 8710,
  8708, 8811, 8448, 8445, 8444, 8443, 8443, 8442, 8441, 8438, 8438, 8438, 
    8438, 8438, 8438, 8650, 8367, 8367, 8367, 8367, 8367, 8367,
  8747, 8846, 8570, 8567, 8565, 8563, 8563, 8562, 8560, 8557, 8557, 8557, 
    8557, 8557, 8557, 8703, 8452, 8452, 8452, 8452, 8452, 8452,
  8643, 8756, 8618, 8621, 8623, 8625, 8628, 8629, 8630, 8633, 8633, 8633, 
    8633, 8633, 8633, 8809, 8764, 8764, 8764, 8764, 8764, 8764,
  8961, 9050, 8605, 8601, 8598, 8596, 8594, 8593, 8591, 8586, 8586, 8586, 
    8586, 8586, 8586, 8775, 8435, 8435, 8435, 8435, 8435, 8435,
  8865, 8958, 8487, 8484, 8482, 8481, 8480, 8480, 8478, 8475, 8475, 8475, 
    8475, 8475, 8475, 8701, 8381, 8381, 8381, 8381, 8381, 8381,
  8530, 8641, 8288, 8287, 8286, 8286, 8286, 8286, 8285, 8284, 8284, 8284, 
    8284, 8284, 8284, 8528, 8253, 8253, 8253, 8253, 8253, 8253,
  8466, 8593, 8534, 8539, 8543, 8545, 8549, 8551, 8553, 8558, 8558, 8558, 
    8558, 8558, 8558, 8757, 8763, 8763, 8763, 8763, 8763, 8763,
  8472, 8599, 8480, 8485, 8489, 8492, 8497, 8499, 8501, 8507, 8507, 8507, 
    8507, 8507, 8507, 8738, 8734, 8734, 8734, 8734, 8734, 8734,
  8448, 8576, 8407, 8413, 8417, 8421, 8425, 8427, 8429, 8436, 8436, 8436, 
    8436, 8436, 8436, 8699, 8678, 8678, 8678, 8678, 8678, 8678,
  8350, 8483, 8313, 8320, 8326, 8329, 8334, 8337, 8339, 8347, 8347, 8347, 
    8347, 8347, 8347, 8638, 8626, 8626, 8626, 8626, 8626, 8626,
  8266, 8401, 8280, 8285, 8289, 8292, 8296, 8298, 8300, 8306, 8306, 8306, 
    8306, 8306, 8306, 8570, 8524, 8524, 8524, 8524, 8524, 8524,
  8207, 8345, 8214, 8219, 8223, 8226, 8230, 8232, 8234, 8239, 8239, 8239, 
    8239, 8239, 8239, 8516, 8448, 8448, 8448, 8448, 8448, 8448,
  8380, 8523, 8153, 8160, 8165, 8169, 8174, 8176, 8178, 8186, 8186, 8186, 
    8186, 8186, 8186, 8626, 8459, 8459, 8459, 8459, 8459, 8459,
  8504, 8640, 8216, 8223, 8228, 8231, 8236, 8238, 8241, 8248, 8248, 8248, 
    8248, 8248, 8248, 8685, 8509, 8509, 8509, 8509, 8509, 8509,
  8606, 8728, 8409, 8413, 8415, 8417, 8419, 8421, 8422, 8425, 8425, 8425, 
    8425, 8425, 8425, 8733, 8560, 8560, 8560, 8560, 8560, 8560,
  8867, 8985, 8895, 8902, 8906, 8909, 8914, 8916, 8918, 8925, 8925, 8925, 
    8925, 8925, 8925, 9124, 9174, 9174, 9174, 9174, 9174, 9174,
  9091, 9196, 9085, 9087, 9088, 9088, 9090, 9090, 9091, 9092, 9092, 9092, 
    9092, 9092, 9092, 9217, 9151, 9151, 9151, 9151, 9151, 9151,
  9292, 9384, 9164, 9168, 9170, 9172, 9175, 9177, 9178, 9182, 9182, 9182, 
    9182, 9182, 9182, 9332, 9335, 9335, 9335, 9335, 9335, 9335,
  9443, 9526, 9230, 9231, 9232, 9233, 9235, 9235, 9236, 9238, 9238, 9238, 
    9238, 9238, 9238, 9373, 9304, 9304, 9304, 9304, 9304, 9304,
  9455, 9547, 9132, 9136, 9139, 9141, 9144, 9145, 9147, 9151, 9151, 9151, 
    9151, 9151, 9151, 9407, 9310, 9310, 9310, 9310, 9310, 9310,
  9434, 9519, 9079, 9088, 9094, 9098, 9103, 9106, 9109, 9118, 9118, 9118, 
    9118, 9118, 9118, 9379, 9436, 9436, 9436, 9436, 9436, 9436,
  9364, 9453, 9050, 9055, 9058, 9060, 9063, 9065, 9066, 9071, 9071, 9071, 
    9071, 9071, 9071, 9308, 9246, 9246, 9246, 9246, 9246, 9246,
  9294, 9388, 9083, 9090, 9094, 9097, 9102, 9104, 9106, 9113, 9113, 9113, 
    9113, 9113, 9113, 9330, 9360, 9360, 9360, 9360, 9360, 9360,
  9209, 9306, 9180, 9185, 9187, 9190, 9193, 9194, 9196, 9200, 9200, 9200, 
    9200, 9200, 9200, 9322, 9367, 9367, 9367, 9367, 9367, 9367,
  8974, 9091, 9085, 9091, 9095, 9098, 9102, 9104, 9107, 9113, 9113, 9113, 
    9113, 9113, 9113, 9264, 9346, 9346, 9346, 9346, 9346, 9346,
  8678, 8816, 8803, 8814, 8822, 8827, 8834, 8837, 8841, 8853, 8853, 8853, 
    8853, 8853, 8853, 9118, 9263, 9263, 9263, 9263, 9263, 9263,
  8334, 8489, 8412, 8429, 8441, 8450, 8460, 8465, 8471, 8490, 8490, 8490, 
    8490, 8490, 8490, 8893, 9135, 9135, 9135, 9135, 9135, 9135,
  8021, 8190, 8049, 8068, 8081, 8091, 8102, 8108, 8115, 8136, 8136, 8136, 
    8136, 8136, 8136, 8628, 8843, 8843, 8843, 8843, 8843, 8843,
  7674, 7852, 7416, 7437, 7451, 7462, 7474, 7482, 7489, 7512, 7512, 7512, 
    7512, 7512, 7512, 8202, 8303, 8303, 8303, 8303, 8303, 8303,
  7206, 7351, 6864, 6881, 6894, 6904, 6913, 6919, 6926, 6946, 6946, 6946, 
    6946, 6946, 6946, 8028, 7824, 7938, 7938, 7938, 7938, 7938,
  6976, 7005, 6156, 6198, 6228, 6251, 6273, 6287, 6302, 6348, 6348, 6348, 
    6348, 6348, 6348, 7345, 7918, 7918, 7918, 7918, 7918, 7918,
  6863, 6893, 6064, 6106, 6136, 6158, 6180, 6194, 6209, 6255, 6255, 6255, 
    6255, 6255, 6255, 7230, 7812, 7811, 7812, 7812, 7811, 7811,
  7146, 7349, 7000, 7019, 7032, 7042, 7053, 7060, 7066, 7087, 7087, 7087, 
    7087, 7087, 7087, 7810, 7796, 7796, 7796, 7796, 7795, 7796,
  7040, 7246, 7669, 7685, 7695, 7703, 7713, 7718, 7723, 7740, 7740, 7740, 
    7740, 7740, 7740, 8057, 8324, 8324, 8324, 8324, 8324, 8324,
  7238, 7440, 8103, 8122, 8135, 8145, 8156, 8162, 8169, 8190, 8190, 8190, 
    8190, 8190, 8190, 8391, 8906, 8905, 8905, 8905, 8905, 8905,
  7550, 7727, 8039, 8051, 8060, 8066, 8074, 8078, 8082, 8096, 8096, 8096, 
    8096, 8096, 8096, 8343, 8569, 8569, 8569, 8569, 8569, 8569,
  7744, 7915, 7811, 7825, 7835, 7843, 7852, 7857, 7862, 7878, 7878, 7878, 
    7878, 7878, 7878, 8329, 8423, 8423, 8423, 8423, 8423, 8423,
  7680, 7856, 7511, 7529, 7542, 7552, 7563, 7569, 7575, 7596, 7596, 7596, 
    7596, 7596, 7596, 8214, 8287, 8287, 8287, 8287, 8287, 8287,
  7281, 7486, 7044, 7068, 7085, 7098, 7112, 7121, 7129, 7156, 7156, 7156, 
    7156, 7156, 7156, 7976, 8072, 8072, 8072, 8072, 8072, 8072,
  7249, 7455, 6999, 7022, 7038, 7050, 7063, 7071, 7079, 7105, 7105, 7105, 
    7105, 7105, 7105, 7923, 7969, 7969, 7969, 7969, 7969, 7969,
  6983, 7155, 6642, 6663, 6678, 6689, 6700, 6707, 6716, 6740, 6740, 6740, 
    6740, 6740, 6740, 7959, 7744, 7866, 7866, 7866, 7866, 7866,
  7151, 7229, 6826, 6859, 6882, 6899, 6916, 6927, 6939, 6975, 6975, 6975, 
    6975, 6975, 6975, 7525, 8182, 8182, 8182, 8182, 8182, 8182,
  7133, 7275, 7150, 7173, 7189, 7201, 7213, 7220, 7229, 7254, 7254, 7254, 
    7254, 7254, 7254, 7595, 8100, 8100, 8100, 8100, 8100, 8100,
  7152, 7402, 7560, 7571, 7579, 7584, 7590, 7593, 7597, 7609, 7609, 7609, 
    7609, 7609, 7609, 7851, 8010, 8010, 8010, 8010, 8010, 8010,
  7282, 7606, 7915, 7917, 7919, 7920, 7921, 7921, 7922, 7925, 7925, 7925, 
    7925, 7925, 7925, 8144, 8000, 8000, 8000, 8000, 8001, 8001,
  7142, 7510, 7958, 7957, 7956, 7955, 7955, 7954, 7953, 7952, 7952, 7952, 
    7952, 7952, 7952, 8116, 7899, 7898, 7898, 7898, 7899, 7899,
  6616, 7041, 7671, 7673, 7674, 7675, 7676, 7676, 7677, 7679, 7679, 7679, 
    7679, 7679, 7679, 7859, 7740, 7740, 7740, 7740, 7740, 7740,
  6216, 6461, 7131, 7159, 7178, 7193, 7207, 7217, 7227, 7258, 7258, 7258, 
    7258, 7258, 7258, 7452, 8253, 8358, 8358, 8358, 8358, 8358,
  5890, 6086, 6834, 6858, 6876, 6889, 6901, 6909, 6919, 6946, 6946, 6946, 
    6946, 6946, 6946, 6963, 7907, 8015, 8015, 8015, 8015, 8015,
  5806, 6037, 6985, 7012, 7032, 7046, 7060, 7069, 7080, 7111, 7111, 7111, 
    7111, 7111, 7111, 7010, 8103, 8208, 8208, 8208, 8208, 8208,
  5874, 6134, 7313, 7342, 7363, 7378, 7393, 7403, 7414, 7446, 7446, 7446, 
    7446, 7446, 7446, 7154, 8404, 8500, 8500, 8500, 8500, 8500,
  8808, 8913, 9000, 8999, 8998, 8998, 8998, 8998, 8997, 8996, 8996, 8996, 
    8996, 8996, 8996, 8998, 8965, 8965, 8965, 8965, 8965, 8965,
  8887, 8988, 9073, 9073, 9073, 9073, 9074, 9074, 9075, 9075, 9075, 9075, 
    9075, 9075, 9075, 9069, 9096, 9096, 9096, 9096, 9096, 9096,
  8851, 8955, 9012, 9014, 9016, 9017, 9019, 9019, 9020, 9023, 9023, 9023, 
    9023, 9023, 9023, 9055, 9110, 9110, 9110, 9110, 9110, 9110,
  8896, 8998, 8985, 8986, 8986, 8986, 8987, 8987, 8988, 8988, 8988, 8988, 
    8988, 8988, 8988, 9039, 9013, 9013, 9013, 9013, 9013, 9013,
  9000, 9097, 9033, 9035, 9036, 9037, 9040, 9040, 9041, 9043, 9043, 9043, 
    9043, 9043, 9043, 9112, 9130, 9130, 9130, 9130, 9130, 9130,
  9023, 9112, 9093, 9095, 9096, 9097, 9099, 9100, 9101, 9103, 9103, 9103, 
    9103, 9103, 9103, 9113, 9190, 9190, 9190, 9190, 9190, 9190,
  8998, 9090, 9065, 9069, 9071, 9072, 9075, 9076, 9077, 9081, 9081, 9081, 
    9081, 9081, 9081, 9112, 9208, 9208, 9208, 9208, 9208, 9208,
  8983, 9077, 9030, 9035, 9039, 9041, 9045, 9047, 9048, 9054, 9054, 9054, 
    9054, 9054, 9054, 9118, 9250, 9250, 9250, 9250, 9250, 9250,
  8987, 9083, 9033, 9038, 9042, 9044, 9048, 9050, 9051, 9057, 9057, 9057, 
    9057, 9057, 9057, 9131, 9259, 9259, 9259, 9259, 9259, 9259,
  8932, 9031, 8940, 8945, 8949, 8952, 8956, 8957, 8959, 8965, 8965, 8965, 
    8965, 8965, 8965, 9074, 9173, 9173, 9173, 9173, 9173, 9173,
  9034, 9129, 9046, 9054, 9059, 9063, 9068, 9070, 9073, 9081, 9081, 9081, 
    9081, 9081, 9081, 9187, 9367, 9367, 9367, 9367, 9367, 9367,
  8953, 9053, 8905, 8912, 8916, 8920, 8924, 8926, 8929, 8936, 8936, 8936, 
    8936, 8936, 8936, 9084, 9187, 9187, 9187, 9187, 9187, 9187,
  8950, 9049, 8894, 8901, 8905, 8909, 8914, 8916, 8919, 8926, 8926, 8926, 
    8926, 8926, 8926, 9080, 9195, 9195, 9195, 9195, 9195, 9195,
  8963, 9063, 8860, 8866, 8871, 8874, 8879, 8881, 8883, 8890, 8890, 8890, 
    8890, 8890, 8890, 9067, 9142, 9142, 9142, 9142, 9142, 9142,
  8990, 9093, 8902, 8903, 8903, 8904, 8906, 8906, 8906, 8908, 8908, 8908, 
    8908, 8908, 8908, 9060, 8960, 8960, 8960, 8960, 8960, 8960,
  9057, 9152, 9002, 9000, 8999, 8998, 8998, 8997, 8996, 8994, 8994, 8994, 
    8994, 8994, 8994, 9075, 8926, 8926, 8926, 8926, 8926, 8926,
  9080, 9168, 8951, 8944, 8939, 8935, 8933, 8930, 8928, 8920, 8920, 8920, 
    8920, 8920, 8920, 8976, 8673, 8673, 8673, 8673, 8673, 8673,
  8991, 9085, 8809, 8806, 8803, 8801, 8800, 8799, 8798, 8794, 8794, 8794, 
    8794, 8794, 8794, 8925, 8668, 8668, 8668, 8668, 8668, 8668,
  8798, 8910, 8669, 8670, 8670, 8671, 8672, 8672, 8672, 8673, 8673, 8673, 
    8673, 8673, 8673, 8885, 8710, 8710, 8710, 8710, 8710, 8710,
  8945, 9046, 8712, 8711, 8710, 8710, 8711, 8710, 8710, 8709, 8709, 8709, 
    8709, 8709, 8709, 8916, 8691, 8691, 8691, 8691, 8691, 8691,
  9164, 9251, 9044, 9037, 9032, 9028, 9025, 9023, 9020, 9012, 9012, 9012, 
    9012, 9012, 9012, 9059, 8749, 8749, 8749, 8749, 8749, 8749,
  9148, 9234, 8981, 8976, 8972, 8969, 8968, 8966, 8964, 8958, 8958, 8958, 
    8958, 8958, 8958, 9039, 8780, 8780, 8780, 8780, 8780, 8780,
  9177, 9262, 9023, 9017, 9014, 9011, 9009, 9007, 9005, 8999, 8999, 8999, 
    8999, 8999, 8999, 9068, 8814, 8814, 8814, 8814, 8814, 8814,
  9069, 9159, 8906, 8902, 8899, 8897, 8895, 8894, 8892, 8887, 8887, 8887, 
    8887, 8887, 8887, 8987, 8735, 8735, 8735, 8735, 8735, 8735,
  8998, 9097, 8803, 8804, 8805, 8805, 8807, 8807, 8808, 8809, 8809, 8809, 
    8809, 8809, 8809, 9003, 8862, 8862, 8862, 8862, 8862, 8862,
  9117, 9216, 8743, 8744, 8744, 8745, 8746, 8746, 8747, 8748, 8748, 8748, 
    8748, 8748, 8748, 9032, 8789, 8789, 8789, 8789, 8789, 8789,
  8995, 9094, 8558, 8557, 8557, 8557, 8558, 8558, 8558, 8558, 8558, 8558, 
    8558, 8558, 8558, 8867, 8560, 8560, 8560, 8560, 8560, 8560,
  8836, 8946, 8394, 8396, 8397, 8398, 8400, 8401, 8401, 8403, 8403, 8403, 
    8403, 8403, 8403, 8772, 8474, 8474, 8474, 8474, 8474, 8474,
  8807, 8920, 8564, 8565, 8565, 8566, 8567, 8567, 8567, 8568, 8568, 8568, 
    8568, 8568, 8568, 8840, 8605, 8605, 8605, 8605, 8605, 8605,
  8702, 8822, 8468, 8470, 8471, 8472, 8474, 8475, 8475, 8477, 8477, 8477, 
    8477, 8477, 8477, 8784, 8555, 8555, 8555, 8555, 8555, 8555,
  8744, 8855, 8376, 8376, 8376, 8377, 8378, 8378, 8378, 8379, 8379, 8379, 
    8379, 8379, 8379, 8707, 8405, 8405, 8405, 8405, 8405, 8405,
  8793, 8904, 8432, 8434, 8435, 8436, 8437, 8438, 8438, 8440, 8440, 8440, 
    8440, 8440, 8440, 8770, 8509, 8509, 8509, 8509, 8509, 8509,
  8911, 9012, 8554, 8553, 8553, 8552, 8553, 8553, 8552, 8552, 8552, 8552, 
    8552, 8552, 8552, 8820, 8536, 8536, 8536, 8536, 8536, 8536,
  8975, 9071, 8628, 8627, 8626, 8625, 8626, 8625, 8625, 8624, 8624, 8624, 
    8624, 8624, 8624, 8860, 8594, 8594, 8594, 8594, 8594, 8594,
  8764, 8870, 8383, 8384, 8385, 8386, 8387, 8388, 8388, 8390, 8390, 8390, 
    8390, 8390, 8390, 8702, 8445, 8445, 8445, 8445, 8445, 8445,
  8633, 8747, 8388, 8390, 8392, 8393, 8395, 8396, 8397, 8400, 8400, 8400, 
    8400, 8400, 8400, 8687, 8500, 8500, 8500, 8500, 8500, 8500,
  8743, 8849, 8414, 8414, 8414, 8415, 8416, 8416, 8416, 8417, 8417, 8417, 
    8417, 8417, 8417, 8699, 8446, 8446, 8446, 8446, 8446, 8446,
  8878, 8977, 8528, 8527, 8527, 8526, 8527, 8526, 8526, 8525, 8525, 8525, 
    8525, 8525, 8525, 8775, 8499, 8499, 8499, 8499, 8499, 8499,
  8848, 8950, 8531, 8530, 8530, 8530, 8531, 8531, 8531, 8531, 8531, 8531, 
    8531, 8531, 8531, 8784, 8535, 8535, 8536, 8536, 8535, 8535,
  8536, 8657, 8524, 8528, 8531, 8533, 8536, 8537, 8539, 8543, 8543, 8543, 
    8543, 8543, 8543, 8750, 8699, 8699, 8699, 8699, 8699, 8699,
  8805, 8905, 8531, 8528, 8526, 8525, 8525, 8524, 8523, 8520, 8520, 8520, 
    8520, 8520, 8520, 8728, 8438, 8438, 8438, 8438, 8438, 8438,
  8697, 8805, 8561, 8558, 8555, 8553, 8553, 8551, 8550, 8546, 8546, 8546, 
    8546, 8546, 8546, 8711, 8425, 8425, 8425, 8425, 8425, 8425,
  8220, 8358, 8361, 8367, 8371, 8375, 8379, 8381, 8384, 8391, 8391, 8391, 
    8391, 8391, 8391, 8606, 8639, 8639, 8639, 8639, 8639, 8639,
  8115, 8258, 8288, 8296, 8301, 8305, 8310, 8313, 8315, 8323, 8323, 8323, 
    8323, 8323, 8323, 8553, 8613, 8613, 8613, 8613, 8613, 8613,
  8390, 8509, 8225, 8224, 8224, 8224, 8225, 8225, 8225, 8224, 8224, 8224, 
    8224, 8224, 8224, 8472, 8227, 8227, 8227, 8227, 8227, 8227,
  8395, 8512, 8213, 8213, 8212, 8212, 8213, 8214, 8213, 8213, 8213, 8213, 
    8213, 8213, 8213, 8454, 8220, 8220, 8220, 8220, 8220, 8220,
  8512, 8622, 8312, 8311, 8311, 8310, 8311, 8311, 8310, 8309, 8309, 8309, 
    8309, 8309, 8309, 8532, 8288, 8288, 8288, 8288, 8288, 8288,
  8438, 8563, 8450, 8456, 8459, 8462, 8466, 8467, 8469, 8475, 8475, 8475, 
    8475, 8475, 8475, 8691, 8678, 8678, 8678, 8678, 8678, 8678,
  8480, 8603, 8466, 8471, 8474, 8476, 8480, 8481, 8483, 8488, 8488, 8488, 
    8488, 8488, 8488, 8705, 8669, 8669, 8669, 8669, 8669, 8669,
  8803, 8901, 8523, 8521, 8520, 8519, 8519, 8518, 8517, 8515, 8515, 8515, 
    8515, 8515, 8515, 8723, 8459, 8459, 8459, 8459, 8459, 8459,
  8602, 8709, 8310, 8311, 8311, 8312, 8313, 8313, 8313, 8314, 8314, 8314, 
    8314, 8314, 8314, 8577, 8344, 8344, 8344, 8344, 8344, 8344,
  8475, 8593, 8253, 8255, 8257, 8258, 8260, 8261, 8262, 8264, 8264, 8264, 
    8264, 8264, 8264, 8549, 8353, 8353, 8353, 8353, 8353, 8353,
  8469, 8593, 8471, 8477, 8480, 8483, 8487, 8489, 8490, 8496, 8496, 8496, 
    8496, 8496, 8496, 8711, 8700, 8700, 8700, 8700, 8700, 8700,
  8445, 8570, 8399, 8403, 8406, 8409, 8412, 8414, 8415, 8420, 8420, 8420, 
    8420, 8420, 8420, 8661, 8597, 8597, 8597, 8597, 8597, 8597,
  8296, 8429, 8270, 8276, 8279, 8282, 8286, 8288, 8290, 8296, 8296, 8296, 
    8296, 8296, 8296, 8570, 8509, 8509, 8509, 8509, 8509, 8509,
  8108, 8248, 7877, 7876, 7875, 7874, 7875, 7875, 7874, 7873, 7873, 7873, 
    7873, 7873, 7873, 8238, 7840, 7840, 7840, 7840, 7840, 7840,
  8131, 8291, 8029, 8036, 8041, 8044, 8049, 8051, 8053, 8061, 8061, 8061, 
    8061, 8061, 8061, 8512, 8318, 8318, 8318, 8318, 8318, 8318,
  7990, 8146, 7910, 7919, 7924, 7928, 7934, 7937, 7939, 7948, 7948, 7948, 
    7948, 7948, 7948, 8369, 8261, 8261, 8261, 8261, 8261, 8261,
  8175, 8322, 8005, 8011, 8016, 8019, 8024, 8026, 8028, 8035, 8035, 8035, 
    8035, 8035, 8035, 8453, 8286, 8286, 8286, 8286, 8286, 8286,
  8555, 8693, 8320, 8326, 8330, 8333, 8337, 8339, 8341, 8347, 8347, 8347, 
    8347, 8347, 8347, 8761, 8566, 8566, 8566, 8566, 8566, 8566,
  8728, 8848, 8629, 8630, 8631, 8632, 8634, 8634, 8634, 8636, 8636, 8636, 
    8636, 8636, 8636, 8871, 8693, 8693, 8693, 8693, 8693, 8693,
  8913, 9025, 8916, 8917, 8919, 8920, 8921, 8922, 8923, 8925, 8925, 8925, 
    8925, 8925, 8925, 9078, 9000, 9000, 9000, 9000, 9000, 9000,
  9261, 9357, 9142, 9148, 9151, 9154, 9157, 9159, 9161, 9166, 9166, 9166, 
    9166, 9166, 9166, 9337, 9362, 9362, 9362, 9362, 9362, 9362,
  9357, 9444, 9161, 9165, 9167, 9169, 9172, 9173, 9175, 9179, 9179, 9179, 
    9179, 9179, 9179, 9339, 9327, 9327, 9327, 9327, 9327, 9327,
  9488, 9570, 9200, 9204, 9207, 9209, 9212, 9214, 9215, 9220, 9220, 9220, 
    9220, 9220, 9220, 9406, 9383, 9383, 9383, 9383, 9383, 9383,
  9415, 9506, 9148, 9154, 9158, 9160, 9164, 9166, 9168, 9175, 9175, 9175, 
    9175, 9175, 9175, 9406, 9398, 9398, 9398, 9398, 9398, 9398,
  9354, 9444, 9177, 9179, 9181, 9183, 9185, 9186, 9187, 9191, 9191, 9191, 
    9191, 9191, 9191, 9351, 9306, 9306, 9306, 9306, 9306, 9306,
  9156, 9263, 9162, 9167, 9170, 9173, 9176, 9177, 9179, 9184, 9184, 9184, 
    9184, 9184, 9184, 9337, 9366, 9366, 9366, 9366, 9366, 9366,
  8790, 8915, 8946, 8954, 8959, 8963, 8968, 8971, 8974, 8982, 8982, 8982, 
    8982, 8982, 8982, 9155, 9282, 9282, 9282, 9282, 9282, 9282,
  8335, 8485, 8484, 8499, 8510, 8518, 8527, 8532, 8537, 8554, 8554, 8554, 
    8554, 8554, 8554, 8883, 9126, 9126, 9126, 9126, 9126, 9126,
  8003, 8171, 7854, 7875, 7890, 7901, 7914, 7921, 7929, 7953, 7953, 7953, 
    7953, 7953, 7953, 8548, 8763, 8763, 8763, 8763, 8763, 8763,
  7925, 8099, 7529, 7551, 7567, 7579, 7591, 7599, 7607, 7632, 7632, 7632, 
    7632, 7632, 7632, 8388, 8468, 8468, 8468, 8468, 8468, 8468,
  7629, 7815, 7260, 7282, 7298, 7309, 7322, 7330, 7338, 7362, 7362, 7362, 
    7362, 7362, 7362, 8154, 8192, 8192, 8192, 8192, 8192, 8192,
  7295, 7495, 7164, 7186, 7202, 7214, 7227, 7236, 7243, 7269, 7269, 7269, 
    7269, 7269, 7269, 7997, 8127, 8127, 8127, 8127, 8127, 8127,
  7055, 7278, 7089, 7111, 7126, 7138, 7151, 7158, 7166, 7190, 7190, 7190, 
    7190, 7190, 7190, 7935, 8018, 8018, 8018, 8018, 8018, 8018,
  6741, 6974, 6786, 6813, 6832, 6846, 6862, 6871, 6881, 6911, 6911, 6911, 
    6911, 6911, 6911, 7719, 7930, 7930, 7930, 7930, 7930, 7930,
  6752, 6912, 6549, 6588, 6615, 6635, 6655, 6668, 6682, 6725, 6725, 6725, 
    6725, 6725, 6725, 7563, 8158, 8158, 8158, 8158, 8158, 8158,
  6879, 7065, 6784, 6821, 6847, 6867, 6886, 6898, 6911, 6952, 6952, 6952, 
    6952, 6952, 6952, 7764, 8324, 8323, 8323, 8324, 8324, 8323,
  6738, 6961, 7372, 7389, 7400, 7410, 7420, 7426, 7432, 7451, 7451, 7451, 
    7451, 7451, 7451, 7844, 8100, 8100, 8100, 8100, 8100, 8100,
  6754, 6979, 7566, 7589, 7605, 7617, 7631, 7639, 7647, 7673, 7673, 7673, 
    7673, 7673, 7673, 8023, 8547, 8547, 8547, 8547, 8547, 8547,
  7119, 7321, 7416, 7433, 7445, 7454, 7464, 7470, 7476, 7495, 7495, 7495, 
    7495, 7495, 7495, 7972, 8144, 8144, 8144, 8144, 8144, 8144,
  7208, 7426, 7125, 7148, 7165, 7178, 7190, 7198, 7208, 7235, 7235, 7235, 
    7235, 7235, 7235, 8312, 8207, 8319, 8319, 8319, 8319, 8319,
  7003, 7187, 6620, 6642, 6658, 6670, 6682, 6690, 6699, 6725, 6725, 6725, 
    6725, 6725, 6725, 8036, 7766, 7891, 7891, 7891, 7891, 7891,
  6809, 6986, 6352, 6375, 6391, 6403, 6415, 6423, 6432, 6459, 6459, 6459, 
    6459, 6459, 6459, 7855, 7559, 7690, 7690, 7690, 7690, 7690,
  6951, 7085, 6644, 6690, 6722, 6746, 6769, 6784, 6800, 6851, 6851, 6851, 
    6851, 6851, 6851, 7764, 8529, 8529, 8529, 8529, 8529, 8529,
  6957, 7076, 6692, 6733, 6762, 6783, 6804, 6818, 6832, 6877, 6877, 6877, 
    6877, 6877, 6877, 7625, 8384, 8384, 8384, 8384, 8384, 8384,
  6933, 7054, 6803, 6833, 6854, 6870, 6885, 6895, 6906, 6939, 6939, 6939, 
    6939, 6939, 6939, 7426, 8041, 8041, 8041, 8041, 8041, 8041,
  7149, 7383, 7422, 7437, 7448, 7456, 7463, 7468, 7473, 7489, 7489, 7489, 
    7489, 7489, 7489, 7857, 8035, 8035, 8035, 8035, 8035, 8035,
  7338, 7636, 7873, 7876, 7879, 7881, 7882, 7883, 7884, 7888, 7888, 7888, 
    7888, 7888, 7888, 8113, 8004, 8004, 8004, 8004, 8004, 8004,
  7354, 7646, 7965, 7960, 7956, 7954, 7951, 7949, 7947, 7941, 7941, 7941, 
    7941, 7941, 7941, 7963, 7742, 7742, 7742, 7742, 7742, 7742,
  7266, 7613, 8053, 8046, 8042, 8038, 8034, 8032, 8029, 8022, 8022, 8022, 
    8022, 8022, 8022, 8072, 7768, 7768, 7768, 7768, 7768, 7768,
  6979, 7401, 7934, 7935, 7936, 7937, 7938, 7938, 7938, 7939, 7939, 7939, 
    7939, 7939, 7939, 8215, 7980, 7980, 7980, 7980, 7981, 7981,
  6263, 6645, 7225, 7232, 7237, 7240, 7244, 7246, 7248, 7256, 7256, 7256, 
    7256, 7256, 7256, 7404, 7509, 7509, 7509, 7509, 7509, 7509,
  5975, 6350, 6964, 6971, 6976, 6980, 6984, 6985, 6988, 6995, 6995, 6995, 
    6995, 6995, 6995, 7084, 7250, 7250, 7250, 7249, 7250, 7250,
  5930, 6180, 7266, 7294, 7314, 7329, 7344, 7353, 7364, 7395, 7395, 7395, 
    7395, 7395, 7395, 7174, 8347, 8444, 8444, 8444, 8444, 8444,
  5584, 6170, 7372, 7361, 7354, 7349, 7343, 7339, 7335, 7322, 7322, 7322, 
    7322, 7322, 7322, 7238, 6912, 6912, 6912, 6912, 6912, 6913,
  8802, 8908, 9031, 9029, 9029, 9028, 9028, 9028, 9027, 9026, 9026, 9026, 
    9026, 9026, 9026, 9009, 8992, 8992, 8992, 8992, 8992, 8992,
  8811, 8912, 9029, 9030, 9031, 9031, 9033, 9033, 9033, 9034, 9034, 9034, 
    9034, 9034, 9034, 9014, 9079, 9079, 9079, 9079, 9079, 9079,
  8816, 8919, 8989, 8989, 8990, 8990, 8991, 8991, 8991, 8992, 8992, 8992, 
    8992, 8992, 8992, 9002, 9018, 9018, 9018, 9018, 9018, 9018,
  8885, 8985, 9052, 9052, 9052, 9052, 9053, 9053, 9053, 9053, 9053, 9053, 
    9053, 9053, 9053, 9051, 9063, 9063, 9063, 9063, 9063, 9063,
  8973, 9065, 9091, 9093, 9095, 9096, 9099, 9099, 9100, 9103, 9103, 9103, 
    9103, 9103, 9103, 9106, 9204, 9204, 9204, 9204, 9204, 9204,
  8963, 9057, 8990, 8992, 8993, 8994, 8996, 8997, 8998, 9000, 9000, 9000, 
    9000, 9000, 9000, 9052, 9083, 9083, 9083, 9083, 9083, 9083,
  9038, 9126, 9103, 9108, 9111, 9114, 9117, 9119, 9121, 9126, 9126, 9126, 
    9126, 9126, 9126, 9151, 9311, 9311, 9311, 9311, 9311, 9311,
  9023, 9115, 9072, 9078, 9082, 9085, 9089, 9090, 9092, 9099, 9099, 9099, 
    9099, 9099, 9099, 9155, 9314, 9314, 9314, 9314, 9314, 9314,
  8979, 9073, 9061, 9066, 9069, 9072, 9075, 9077, 9078, 9084, 9084, 9084, 
    9084, 9084, 9084, 9130, 9269, 9269, 9269, 9269, 9269, 9269,
  9007, 9102, 9077, 9085, 9091, 9095, 9100, 9102, 9105, 9114, 9114, 9114, 
    9114, 9114, 9114, 9188, 9414, 9414, 9414, 9414, 9414, 9414,
  8980, 9076, 9028, 9035, 9040, 9044, 9049, 9051, 9054, 9062, 9062, 9062, 
    9062, 9062, 9062, 9150, 9336, 9336, 9336, 9336, 9336, 9336,
  8936, 9033, 8969, 8975, 8980, 8983, 8988, 8990, 8992, 9000, 9000, 9000, 
    9000, 9000, 9000, 9093, 9252, 9252, 9252, 9252, 9252, 9252,
  8895, 8991, 8881, 8886, 8890, 8893, 8897, 8899, 8901, 8907, 8907, 8907, 
    8907, 8907, 8907, 9015, 9126, 9126, 9126, 9126, 9126, 9126,
  9048, 9145, 9001, 9007, 9011, 9014, 9018, 9020, 9022, 9028, 9028, 9028, 
    9028, 9028, 9028, 9158, 9245, 9245, 9245, 9245, 9245, 9245,
  9067, 9164, 9041, 9039, 9038, 9037, 9037, 9036, 9036, 9034, 9034, 9034, 
    9034, 9034, 9034, 9114, 8980, 8980, 8980, 8980, 8980, 8980,
  9085, 9176, 8998, 8994, 8992, 8991, 8990, 8989, 8988, 8984, 8984, 8984, 
    8984, 8984, 8984, 9056, 8879, 8879, 8879, 8879, 8879, 8879,
  9053, 9143, 8845, 8842, 8839, 8837, 8836, 8835, 8834, 8830, 8830, 8830, 
    8830, 8830, 8830, 8956, 8706, 8706, 8706, 8706, 8706, 8706,
  8683, 8802, 8603, 8605, 8607, 8608, 8610, 8610, 8611, 8613, 8613, 8613, 
    8613, 8613, 8613, 8836, 8694, 8694, 8694, 8694, 8694, 8694,
  8587, 8714, 8495, 8497, 8499, 8501, 8503, 8504, 8505, 8509, 8509, 8509, 
    8509, 8509, 8509, 8781, 8625, 8625, 8625, 8625, 8625, 8625,
  8988, 9085, 8789, 8788, 8787, 8786, 8786, 8786, 8785, 8784, 8784, 8784, 
    8784, 8784, 8784, 8948, 8742, 8742, 8742, 8742, 8742, 8742,
  9099, 9189, 9016, 9009, 9005, 9002, 8999, 8997, 8995, 8988, 8988, 8988, 
    8988, 8988, 8988, 9032, 8765, 8765, 8765, 8765, 8765, 8765,
  9091, 9179, 8948, 8943, 8939, 8936, 8934, 8932, 8930, 8923, 8923, 8923, 
    8923, 8923, 8923, 8996, 8722, 8722, 8722, 8722, 8722, 8722,
  9106, 9193, 8964, 8958, 8953, 8949, 8947, 8944, 8942, 8934, 8934, 8934, 
    8934, 8934, 8934, 8994, 8692, 8693, 8693, 8693, 8693, 8693,
  9070, 9161, 8900, 8894, 8890, 8888, 8886, 8884, 8882, 8876, 8876, 8876, 
    8876, 8876, 8876, 8976, 8683, 8683, 8683, 8683, 8683, 8683,
  9098, 9192, 8777, 8775, 8773, 8772, 8772, 8771, 8770, 8768, 8768, 8768, 
    8768, 8768, 8768, 8982, 8690, 8690, 8691, 8691, 8690, 8690,
  9100, 9199, 8570, 8571, 8571, 8572, 8573, 8574, 8574, 8575, 8575, 8575, 
    8575, 8575, 8575, 8936, 8620, 8620, 8620, 8620, 8620, 8620,
  8998, 9098, 8561, 8561, 8561, 8560, 8561, 8561, 8561, 8561, 8561, 8561, 
    8561, 8561, 8561, 8871, 8557, 8557, 8557, 8557, 8557, 8557,
  8844, 8953, 8545, 8546, 8546, 8547, 8548, 8549, 8549, 8550, 8550, 8550, 
    8550, 8550, 8550, 8834, 8590, 8590, 8590, 8590, 8590, 8590,
  8883, 8994, 8602, 8603, 8604, 8605, 8606, 8607, 8607, 8608, 8608, 8608, 
    8608, 8608, 8608, 8897, 8658, 8658, 8658, 8658, 8658, 8658,
  8959, 9068, 8713, 8714, 8714, 8714, 8715, 8716, 8716, 8716, 8716, 8716, 
    8716, 8716, 8716, 8973, 8745, 8745, 8745, 8745, 8745, 8745,
  8971, 9073, 8664, 8663, 8663, 8663, 8663, 8663, 8663, 8663, 8663, 8663, 
    8663, 8663, 8663, 8916, 8657, 8657, 8657, 8657, 8657, 8657,
  8956, 9057, 8589, 8588, 8588, 8588, 8588, 8588, 8588, 8587, 8587, 8587, 
    8587, 8587, 8587, 8864, 8578, 8578, 8578, 8578, 8578, 8578,
  8719, 8832, 8688, 8690, 8692, 8694, 8697, 8698, 8699, 8702, 8702, 8702, 
    8702, 8702, 8702, 8879, 8822, 8822, 8822, 8822, 8822, 8822,
  8662, 8778, 8663, 8667, 8670, 8671, 8674, 8676, 8677, 8681, 8681, 8681, 
    8681, 8681, 8681, 8858, 8826, 8826, 8826, 8826, 8826, 8826,
  8600, 8719, 8643, 8647, 8649, 8651, 8654, 8656, 8657, 8662, 8662, 8662, 
    8662, 8662, 8662, 8833, 8818, 8818, 8818, 8818, 8818, 8818,
  8547, 8669, 8612, 8615, 8618, 8620, 8623, 8624, 8625, 8630, 8630, 8630, 
    8630, 8630, 8630, 8801, 8778, 8778, 8778, 8778, 8778, 8778,
  8519, 8643, 8590, 8594, 8597, 8599, 8602, 8603, 8604, 8609, 8609, 8609, 
    8609, 8609, 8609, 8784, 8763, 8763, 8763, 8763, 8763, 8763,
  8653, 8768, 8655, 8658, 8660, 8661, 8664, 8665, 8666, 8669, 8669, 8669, 
    8669, 8669, 8669, 8831, 8784, 8784, 8783, 8783, 8784, 8784,
  8581, 8699, 8615, 8619, 8622, 8624, 8627, 8628, 8630, 8634, 8634, 8634, 
    8634, 8634, 8634, 8804, 8789, 8789, 8789, 8789, 8789, 8789,
  8508, 8631, 8537, 8541, 8545, 8547, 8551, 8552, 8554, 8559, 8559, 8559, 
    8559, 8559, 8559, 8758, 8743, 8743, 8743, 8743, 8743, 8743,
  8496, 8618, 8471, 8476, 8478, 8481, 8484, 8485, 8487, 8491, 8491, 8491, 
    8491, 8491, 8491, 8709, 8657, 8657, 8657, 8657, 8657, 8657,
  8507, 8622, 8324, 8323, 8322, 8322, 8322, 8322, 8322, 8321, 8321, 8321, 
    8321, 8321, 8321, 8554, 8301, 8301, 8301, 8301, 8301, 8301,
  8168, 8309, 8294, 8301, 8306, 8310, 8315, 8318, 8320, 8328, 8328, 8328, 
    8328, 8328, 8328, 8570, 8610, 8610, 8610, 8610, 8610, 8610,
  8166, 8308, 8277, 8283, 8288, 8292, 8297, 8299, 8301, 8309, 8309, 8309, 
    8309, 8309, 8309, 8557, 8575, 8575, 8575, 8575, 8575, 8575,
  8394, 8539, 8309, 8298, 8291, 8286, 8281, 8278, 8274, 8263, 8263, 8263, 
    8263, 8263, 8263, 8535, 7892, 7892, 7892, 7892, 7892, 7892,
  8175, 8304, 8121, 8124, 8125, 8127, 8129, 8130, 8131, 8134, 8134, 8134, 
    8134, 8134, 8134, 8379, 8239, 8239, 8239, 8239, 8239, 8239,
  8169, 8309, 8268, 8276, 8281, 8285, 8290, 8293, 8296, 8304, 8304, 8304, 
    8304, 8304, 8304, 8561, 8600, 8600, 8600, 8600, 8600, 8600,
  8183, 8324, 8320, 8327, 8332, 8336, 8341, 8344, 8346, 8355, 8355, 8355, 
    8355, 8355, 8355, 8592, 8643, 8643, 8643, 8643, 8643, 8643,
  8213, 8342, 8147, 8149, 8150, 8151, 8153, 8153, 8154, 8156, 8156, 8156, 
    8156, 8156, 8156, 8405, 8228, 8228, 8228, 8228, 8228, 8228,
  8371, 8500, 8450, 8455, 8459, 8462, 8465, 8467, 8469, 8475, 8475, 8475, 
    8475, 8475, 8475, 8679, 8687, 8687, 8687, 8687, 8687, 8687,
  8288, 8422, 8361, 8367, 8371, 8375, 8379, 8381, 8383, 8390, 8390, 8390, 
    8390, 8390, 8390, 8621, 8635, 8635, 8635, 8635, 8635, 8635,
  8368, 8497, 8425, 8430, 8434, 8437, 8441, 8443, 8445, 8451, 8451, 8451, 
    8451, 8451, 8451, 8662, 8670, 8670, 8670, 8670, 8670, 8670,
  8483, 8597, 8223, 8221, 8220, 8219, 8219, 8219, 8218, 8216, 8216, 8216, 
    8216, 8216, 8216, 8477, 8164, 8164, 8164, 8164, 8164, 8164,
  8189, 8327, 8225, 8230, 8234, 8237, 8241, 8243, 8245, 8251, 8251, 8251, 
    8251, 8251, 8251, 8513, 8465, 8465, 8465, 8465, 8465, 8465,
  8008, 8157, 8114, 8121, 8125, 8129, 8133, 8136, 8138, 8145, 8145, 8145, 
    8145, 8145, 8145, 8424, 8400, 8400, 8400, 8400, 8400, 8400,
  7978, 8139, 7999, 8004, 8006, 8009, 8012, 8014, 8015, 8020, 8020, 8020, 
    8020, 8020, 8020, 8393, 8188, 8188, 8188, 8188, 8188, 8188,
  7826, 7999, 7675, 7688, 7697, 7704, 7712, 7716, 7721, 7735, 7735, 7735, 
    7735, 7735, 7735, 8302, 8230, 8230, 8230, 8230, 8230, 8230,
  7813, 7980, 7713, 7722, 7728, 7733, 7739, 7743, 7746, 7756, 7756, 7756, 
    7756, 7756, 7756, 8239, 8110, 8110, 8110, 8110, 8110, 8110,
  7925, 8087, 7772, 7781, 7786, 7791, 7796, 7799, 7802, 7811, 7811, 7811, 
    7811, 7811, 7811, 8299, 8132, 8132, 8132, 8132, 8132, 8132,
  8180, 8326, 7975, 7980, 7984, 7987, 7991, 7993, 7994, 8000, 8000, 8000, 
    8000, 8000, 8000, 8427, 8212, 8212, 8212, 8212, 8212, 8212,
  8509, 8637, 8369, 8370, 8370, 8371, 8372, 8372, 8373, 8374, 8374, 8374, 
    8374, 8374, 8374, 8660, 8415, 8415, 8415, 8415, 8415, 8415,
  8700, 8825, 8846, 8853, 8858, 8862, 8867, 8869, 8872, 8880, 8880, 8880, 
    8880, 8880, 8880, 9055, 9164, 9164, 9164, 9164, 9164, 9164,
  8956, 9069, 9032, 9039, 9044, 9047, 9052, 9054, 9057, 9065, 9065, 9065, 
    9065, 9065, 9065, 9219, 9333, 9333, 9333, 9333, 9333, 9333,
  9228, 9328, 9207, 9214, 9219, 9223, 9227, 9230, 9232, 9240, 9240, 9240, 
    9240, 9240, 9240, 9391, 9515, 9515, 9515, 9515, 9514, 9515,
  9292, 9385, 9196, 9199, 9202, 9203, 9206, 9207, 9208, 9211, 9211, 9211, 
    9211, 9211, 9211, 9340, 9333, 9333, 9333, 9333, 9333, 9333,
  9165, 9267, 9137, 9139, 9140, 9141, 9143, 9144, 9144, 9146, 9146, 9146, 
    9146, 9146, 9146, 9275, 9227, 9227, 9227, 9227, 9227, 9227,
  8933, 9048, 9015, 9022, 9027, 9030, 9035, 9037, 9039, 9047, 9047, 9047, 
    9047, 9047, 9047, 9204, 9307, 9307, 9307, 9307, 9307, 9307,
  8697, 8833, 8841, 8857, 8867, 8875, 8885, 8890, 8895, 8913, 8913, 8913, 
    8913, 8913, 8913, 9187, 9497, 9497, 9497, 9497, 9497, 9497,
  8178, 8343, 8199, 8224, 8241, 8253, 8267, 8276, 8284, 8311, 8311, 8311, 
    8311, 8311, 8311, 8830, 9228, 9228, 9228, 9228, 9228, 9228,
  7779, 7951, 7576, 7601, 7619, 7633, 7647, 7656, 7665, 7694, 7694, 7694, 
    7694, 7694, 7694, 8354, 8661, 8661, 8661, 8661, 8661, 8661,
  7791, 7978, 7270, 7292, 7307, 7319, 7332, 7340, 7347, 7372, 7372, 7372, 
    7372, 7372, 7372, 8249, 8205, 8205, 8205, 8205, 8205, 8205,
  7261, 7401, 6696, 6714, 6726, 6736, 6745, 6751, 6758, 6779, 6779, 6779, 
    6779, 6779, 6779, 8090, 7702, 7822, 7822, 7822, 7822, 7822,
  6984, 7157, 6575, 6596, 6612, 6624, 6635, 6642, 6651, 6676, 6676, 6676, 
    6676, 6676, 6676, 7979, 7705, 7830, 7830, 7830, 7830, 7830,
  6835, 7068, 6642, 6668, 6687, 6701, 6715, 6725, 6734, 6763, 6763, 6763, 
    6763, 6763, 6763, 7692, 7748, 7748, 7748, 7748, 7748, 7748,
  6414, 6658, 6998, 7014, 7026, 7036, 7046, 7052, 7058, 7077, 7077, 7077, 
    7077, 7077, 7077, 7594, 7729, 7729, 7728, 7728, 7729, 7729,
  5966, 6228, 6510, 6543, 6566, 6584, 6603, 6615, 6626, 6663, 6663, 6663, 
    6663, 6663, 6663, 7370, 7921, 7921, 7921, 7921, 7921, 7921,
  6447, 6703, 6449, 6479, 6500, 6516, 6533, 6544, 6554, 6588, 6588, 6588, 
    6588, 6588, 6588, 7539, 7720, 7720, 7720, 7720, 7720, 7720,
  6412, 6595, 6332, 6356, 6373, 6386, 6398, 6406, 6416, 6443, 6443, 6443, 
    6443, 6443, 6443, 7487, 7542, 7670, 7670, 7670, 7670, 7670,
  6437, 6682, 6780, 6804, 6821, 6833, 6847, 6855, 6864, 6890, 6890, 6890, 
    6890, 6890, 6890, 7574, 7789, 7789, 7789, 7789, 7789, 7789,
  6288, 6537, 6657, 6686, 6707, 6723, 6739, 6750, 6760, 6793, 6793, 6793, 
    6793, 6793, 6793, 7516, 7906, 7906, 7906, 7906, 7906, 7906,
  6841, 7071, 6729, 6752, 6768, 6780, 6793, 6802, 6810, 6835, 6835, 6835, 
    6835, 6835, 6835, 7693, 7708, 7708, 7708, 7708, 7708, 7708,
  6615, 6811, 6249, 6274, 6292, 6305, 6318, 6327, 6337, 6366, 6366, 6366, 
    6366, 6366, 6366, 7762, 7537, 7672, 7672, 7672, 7672, 7672,
  6623, 6740, 6092, 6144, 6180, 6207, 6234, 6252, 6270, 6327, 6327, 6327, 
    6327, 6327, 6327, 7483, 8243, 8243, 8243, 8243, 8243, 8243,
  6566, 6681, 6189, 6242, 6279, 6306, 6334, 6351, 6370, 6428, 6428, 6428, 
    6428, 6428, 6428, 7413, 8375, 8375, 8375, 8375, 8375, 8375,
  6600, 6724, 6362, 6411, 6445, 6470, 6495, 6511, 6528, 6581, 6581, 6581, 
    6581, 6581, 6581, 7404, 8367, 8366, 8366, 8367, 8367, 8366,
  6687, 6863, 6683, 6718, 6743, 6761, 6779, 6791, 6804, 6842, 6842, 6842, 
    6842, 6842, 6842, 7486, 8141, 8141, 8141, 8141, 8141, 8141,
  6895, 7148, 7235, 7256, 7270, 7281, 7291, 7298, 7305, 7328, 7328, 7328, 
    7328, 7328, 7328, 7765, 8086, 8086, 8086, 8086, 8086, 8086,
  7188, 7449, 7590, 7601, 7609, 7614, 7619, 7622, 7626, 7637, 7637, 7637, 
    7637, 7637, 7637, 7932, 8019, 8019, 8019, 8019, 8019, 8019,
  7574, 7861, 8078, 8077, 8077, 8077, 8077, 8076, 8076, 8075, 8075, 8075, 
    8075, 8075, 8075, 8248, 8048, 8048, 8048, 8048, 8048, 8049,
  7749, 8037, 8264, 8258, 8254, 8251, 8248, 8245, 8243, 8237, 8237, 8237, 
    8237, 8237, 8237, 8344, 8011, 8011, 8011, 8011, 8012, 8012,
  7592, 7901, 8200, 8197, 8194, 8192, 8190, 8188, 8187, 8183, 8183, 8183, 
    8183, 8183, 8183, 8303, 8039, 8039, 8039, 8039, 8039, 8039,
  7113, 7511, 8024, 8021, 8020, 8018, 8016, 8015, 8014, 8010, 8010, 8010, 
    8010, 8010, 8010, 8183, 7896, 7896, 7896, 7896, 7896, 7896,
  6567, 6941, 7499, 7501, 7503, 7504, 7504, 7505, 7505, 7507, 7507, 7507, 
    7507, 7507, 7507, 7602, 7570, 7570, 7570, 7570, 7570, 7570,
  6158, 6524, 7124, 7128, 7131, 7133, 7135, 7136, 7137, 7141, 7141, 7141, 
    7141, 7141, 7141, 7180, 7274, 7274, 7274, 7274, 7274, 7274,
  5890, 6418, 7360, 7359, 7359, 7358, 7357, 7357, 7356, 7355, 7355, 7355, 
    7355, 7355, 7355, 7486, 7309, 7309, 7309, 7309, 7309, 7310,
  5652, 6254, 7482, 7471, 7463, 7457, 7451, 7446, 7442, 7429, 7429, 7429, 
    7429, 7429, 7429, 7360, 6991, 6991, 6991, 6991, 6991, 6991,
  8806, 8913, 9062, 9061, 9061, 9061, 9061, 9061, 9061, 9061, 9061, 9061, 
    9061, 9061, 9061, 9043, 9056, 9056, 9056, 9056, 9056, 9056,
  8810, 8917, 8986, 8988, 8989, 8990, 8992, 8993, 8993, 8995, 8995, 8995, 
    8995, 8995, 8995, 9032, 9075, 9075, 9075, 9075, 9075, 9075,
  8870, 8973, 9071, 9070, 9069, 9069, 9069, 9069, 9069, 9068, 9068, 9068, 
    9068, 9068, 9068, 9057, 9046, 9046, 9046, 9046, 9046, 9046,
  8921, 9028, 9072, 9069, 9067, 9065, 9064, 9063, 9062, 9059, 9059, 9059, 
    9059, 9059, 9059, 9082, 8953, 8953, 8953, 8953, 8953, 8953,
  9007, 9108, 9086, 9086, 9085, 9085, 9086, 9085, 9085, 9084, 9084, 9084, 
    9084, 9084, 9084, 9129, 9070, 9070, 9070, 9070, 9070, 9070,
  8958, 9051, 9044, 9047, 9049, 9051, 9053, 9054, 9055, 9059, 9059, 9059, 
    9059, 9059, 9059, 9087, 9182, 9182, 9182, 9182, 9182, 9182,
  9004, 9098, 9060, 9064, 9067, 9068, 9071, 9073, 9074, 9078, 9078, 9078, 
    9078, 9078, 9078, 9130, 9228, 9228, 9228, 9228, 9228, 9228,
  8973, 9067, 9009, 9014, 9018, 9021, 9025, 9027, 9029, 9035, 9035, 9035, 
    9035, 9035, 9035, 9107, 9246, 9246, 9246, 9246, 9246, 9246,
  9001, 9102, 9076, 9083, 9088, 9091, 9096, 9098, 9101, 9108, 9108, 9108, 
    9108, 9108, 9108, 9207, 9371, 9371, 9371, 9371, 9371, 9371,
  8963, 9065, 9003, 9011, 9016, 9020, 9025, 9027, 9030, 9038, 9038, 9038, 
    9038, 9038, 9038, 9160, 9330, 9330, 9330, 9330, 9330, 9330,
  8926, 9027, 8949, 8957, 8962, 8966, 8971, 8973, 8976, 8985, 8985, 8985, 
    8985, 8985, 8985, 9112, 9281, 9281, 9281, 9281, 9281, 9281,
  8924, 9031, 8913, 8917, 8920, 8922, 8925, 8927, 8928, 8933, 8933, 8933, 
    8933, 8933, 8933, 9082, 9092, 9092, 9092, 9092, 9092, 9092,
  8922, 9026, 8897, 8902, 8905, 8908, 8911, 8913, 8915, 8920, 8920, 8920, 
    8920, 8920, 8920, 9068, 9108, 9108, 9108, 9108, 9108, 9108,
  9026, 9129, 8919, 8920, 8920, 8920, 8922, 8922, 8922, 8922, 8922, 8922, 
    8922, 8922, 8922, 9084, 8949, 8949, 8949, 8949, 8949, 8949,
  9022, 9120, 9005, 9004, 9003, 9003, 9003, 9003, 9002, 9001, 9001, 9001, 
    9001, 9001, 9001, 9085, 8972, 8972, 8972, 8972, 8972, 8972,
  9104, 9194, 9030, 9027, 9024, 9023, 9022, 9021, 9020, 9017, 9017, 9017, 
    9017, 9017, 9017, 9080, 8914, 8914, 8914, 8914, 8914, 8914,
  9245, 9315, 9045, 9034, 9026, 9020, 9015, 9011, 9007, 8995, 8995, 8995, 
    8995, 8995, 8995, 8978, 8587, 8587, 8587, 8587, 8587, 8587,
  8613, 8735, 8518, 8521, 8523, 8524, 8526, 8527, 8528, 8530, 8530, 8530, 
    8530, 8530, 8530, 8779, 8630, 8630, 8630, 8630, 8630, 8630,
  8832, 8937, 8647, 8645, 8643, 8642, 8641, 8640, 8639, 8637, 8637, 8637, 
    8637, 8637, 8637, 8825, 8552, 8552, 8552, 8552, 8552, 8552,
  8965, 9062, 8828, 8823, 8819, 8817, 8815, 8813, 8811, 8805, 8805, 8805, 
    8805, 8805, 8805, 8916, 8619, 8619, 8619, 8619, 8619, 8619,
  8987, 9084, 8821, 8815, 8811, 8808, 8806, 8804, 8802, 8796, 8796, 8796, 
    8796, 8796, 8796, 8918, 8597, 8597, 8597, 8597, 8597, 8597,
  8996, 9091, 8914, 8911, 8908, 8907, 8906, 8904, 8903, 8899, 8899, 8899, 
    8899, 8899, 8899, 8984, 8781, 8781, 8781, 8781, 8781, 8781,
  9009, 9107, 8921, 8921, 8920, 8920, 8921, 8920, 8920, 8919, 8919, 8919, 
    8919, 8919, 8919, 9039, 8907, 8907, 8907, 8907, 8907, 8907,
  9033, 9129, 8870, 8869, 8868, 8867, 8867, 8867, 8867, 8865, 8865, 8865, 
    8865, 8865, 8865, 9011, 8832, 8832, 8832, 8832, 8832, 8832,
  9205, 9295, 8877, 8874, 8872, 8870, 8870, 8869, 8868, 8864, 8864, 8864, 
    8864, 8864, 8864, 9061, 8766, 8766, 8766, 8766, 8766, 8766,
  9139, 9234, 8764, 8762, 8761, 8760, 8761, 8760, 8760, 8758, 8758, 8758, 
    8758, 8758, 8758, 9009, 8715, 8715, 8715, 8715, 8715, 8715,
  8958, 9061, 8660, 8660, 8660, 8660, 8661, 8661, 8661, 8661, 8661, 8661, 
    8661, 8661, 8661, 8917, 8671, 8671, 8671, 8671, 8671, 8671,
  9042, 9140, 8788, 8787, 8785, 8784, 8784, 8784, 8783, 8781, 8781, 8781, 
    8781, 8781, 8781, 8982, 8728, 8728, 8728, 8728, 8728, 8728,
  9194, 9287, 9031, 9028, 9026, 9024, 9023, 9022, 9021, 9017, 9017, 9017, 
    9017, 9017, 9017, 9139, 8909, 8909, 8909, 8909, 8909, 8909,
  9271, 9356, 9052, 9047, 9044, 9041, 9040, 9038, 9036, 9031, 9031, 9031, 
    9031, 9031, 9031, 9137, 8860, 8860, 8860, 8860, 8860, 8860,
  9070, 9168, 8737, 8737, 8737, 8736, 8737, 8737, 8737, 8736, 8736, 8736, 
    8736, 8736, 8736, 8986, 8733, 8733, 8733, 8733, 8733, 8733,
  8716, 8832, 8482, 8484, 8486, 8487, 8489, 8490, 8491, 8494, 8494, 8494, 
    8494, 8494, 8494, 8783, 8596, 8596, 8596, 8596, 8596, 8596,
  8729, 8844, 8733, 8736, 8738, 8739, 8742, 8742, 8744, 8747, 8747, 8747, 
    8747, 8747, 8747, 8913, 8863, 8863, 8863, 8863, 8863, 8863,
  8641, 8761, 8641, 8645, 8648, 8650, 8653, 8654, 8656, 8660, 8660, 8660, 
    8660, 8660, 8660, 8856, 8818, 8818, 8818, 8818, 8818, 8818,
  8591, 8713, 8617, 8622, 8625, 8627, 8631, 8632, 8634, 8639, 8639, 8639, 
    8639, 8639, 8639, 8836, 8815, 8815, 8815, 8815, 8815, 8815,
  8505, 8630, 8555, 8560, 8563, 8565, 8569, 8570, 8572, 8577, 8577, 8577, 
    8577, 8577, 8577, 8778, 8760, 8760, 8760, 8760, 8760, 8760,
  8515, 8639, 8544, 8549, 8552, 8554, 8558, 8559, 8561, 8566, 8566, 8566, 
    8566, 8566, 8566, 8772, 8753, 8753, 8753, 8753, 8753, 8753,
  8425, 8553, 8549, 8553, 8556, 8559, 8562, 8564, 8565, 8570, 8570, 8570, 
    8570, 8570, 8570, 8743, 8746, 8746, 8746, 8746, 8746, 8746,
  8065, 8208, 8023, 8028, 8032, 8035, 8039, 8041, 8043, 8049, 8049, 8049, 
    8049, 8049, 8049, 8374, 8270, 8270, 8270, 8270, 8270, 8270,
  8701, 8807, 8455, 8452, 8450, 8449, 8448, 8447, 8446, 8443, 8443, 8443, 
    8443, 8443, 8443, 8663, 8355, 8355, 8355, 8355, 8355, 8355,
  8658, 8767, 8472, 8466, 8463, 8460, 8458, 8456, 8454, 8448, 8448, 8448, 
    8448, 8448, 8448, 8631, 8259, 8259, 8259, 8259, 8259, 8259,
  8230, 8368, 8346, 8353, 8357, 8360, 8364, 8367, 8369, 8376, 8376, 8376, 
    8376, 8376, 8376, 8605, 8618, 8618, 8618, 8618, 8618, 8618,
  8071, 8219, 8259, 8267, 8273, 8277, 8283, 8286, 8288, 8298, 8298, 8298, 
    8298, 8298, 8298, 8544, 8620, 8620, 8620, 8620, 8620, 8620,
  8048, 8197, 8163, 8172, 8179, 8184, 8189, 8193, 8196, 8206, 8206, 8206, 
    8206, 8206, 8206, 8502, 8558, 8558, 8558, 8558, 8558, 8558,
  8002, 8153, 8113, 8123, 8130, 8135, 8141, 8145, 8148, 8159, 8159, 8159, 
    8159, 8159, 8159, 8472, 8540, 8540, 8540, 8540, 8540, 8540,
  7993, 8144, 8131, 8140, 8146, 8151, 8157, 8160, 8163, 8173, 8173, 8173, 
    8173, 8173, 8173, 8465, 8519, 8519, 8519, 8519, 8519, 8519,
  8081, 8227, 8197, 8206, 8212, 8216, 8222, 8225, 8228, 8237, 8237, 8237, 
    8237, 8237, 8237, 8512, 8564, 8564, 8564, 8564, 8564, 8564,
  8176, 8317, 8233, 8242, 8248, 8253, 8259, 8262, 8265, 8275, 8275, 8275, 
    8275, 8275, 8275, 8562, 8617, 8617, 8617, 8617, 8617, 8617,
  8302, 8434, 8344, 8349, 8353, 8356, 8361, 8363, 8365, 8371, 8371, 8371, 
    8371, 8371, 8371, 8611, 8598, 8598, 8598, 8598, 8598, 8598,
  8363, 8484, 8239, 8238, 8238, 8238, 8239, 8239, 8239, 8239, 8239, 8239, 
    8239, 8239, 8239, 8470, 8243, 8243, 8243, 8243, 8243, 8243,
  8275, 8398, 8145, 8147, 8148, 8149, 8150, 8151, 8151, 8153, 8153, 8153, 
    8153, 8153, 8153, 8405, 8220, 8220, 8220, 8220, 8220, 8220,
  8469, 8582, 8313, 8312, 8311, 8311, 8311, 8311, 8311, 8310, 8310, 8310, 
    8310, 8310, 8310, 8520, 8293, 8293, 8293, 8293, 8293, 8293,
  8243, 8366, 8031, 8029, 8028, 8026, 8026, 8026, 8025, 8022, 8022, 8022, 
    8022, 8022, 8022, 8296, 7950, 7950, 7950, 7950, 7950, 7950,
  8068, 8206, 7873, 7873, 7873, 7873, 7874, 7875, 7874, 7874, 7874, 7874, 
    7874, 7874, 7874, 8221, 7888, 7888, 7888, 7888, 7888, 7888,
  8042, 8207, 8048, 8054, 8058, 8062, 8066, 8068, 8070, 8077, 8077, 8077, 
    8077, 8077, 8077, 8486, 8314, 8314, 8314, 8314, 8314, 8314,
  7680, 7855, 7575, 7587, 7596, 7602, 7610, 7614, 7619, 7632, 7632, 7632, 
    7632, 7632, 7632, 8173, 8102, 8102, 8102, 8102, 8102, 8102,
  7703, 7884, 7396, 7414, 7426, 7436, 7446, 7453, 7459, 7479, 7479, 7479, 
    7479, 7479, 7479, 8190, 8151, 8151, 8151, 8151, 8151, 8151,
  7664, 7839, 7525, 7535, 7542, 7547, 7554, 7557, 7561, 7572, 7572, 7572, 
    7572, 7572, 7572, 8118, 7956, 7956, 7956, 7956, 7956, 7956,
  7688, 7864, 7525, 7541, 7553, 7561, 7571, 7577, 7583, 7601, 7601, 7601, 
    7601, 7601, 7601, 8203, 8224, 8224, 8224, 8224, 8224, 8224,
  7912, 8083, 7697, 7711, 7722, 7730, 7738, 7744, 7749, 7765, 7765, 7765, 
    7765, 7765, 7765, 8366, 8322, 8322, 8322, 8322, 8322, 8322,
  8113, 8264, 8004, 8009, 8013, 8016, 8021, 8023, 8025, 8031, 8031, 8031, 
    8031, 8031, 8031, 8435, 8257, 8257, 8257, 8257, 8257, 8257,
  8290, 8441, 8539, 8549, 8556, 8562, 8568, 8572, 8576, 8588, 8588, 8588, 
    8588, 8588, 8588, 8842, 8991, 8991, 8991, 8991, 8991, 8991,
  8508, 8649, 8858, 8864, 8868, 8872, 8876, 8878, 8880, 8888, 8888, 8888, 
    8888, 8888, 8888, 9023, 9135, 9135, 9135, 9135, 9135, 9135,
  8682, 8812, 8926, 8931, 8935, 8938, 8941, 8943, 8945, 8951, 8951, 8951, 
    8951, 8951, 8951, 9080, 9150, 9150, 9150, 9150, 9150, 9150,
  8633, 8762, 8779, 8781, 8783, 8784, 8786, 8787, 8788, 8791, 8791, 8791, 
    8791, 8791, 8791, 8952, 8896, 8896, 8896, 8896, 8896, 8896,
  8596, 8734, 8843, 8850, 8856, 8860, 8865, 8868, 8870, 8879, 8879, 8879, 
    8879, 8879, 8879, 9063, 9181, 9181, 9181, 9181, 9181, 9181,
  8327, 8481, 8561, 8580, 8594, 8604, 8615, 8622, 8628, 8650, 8650, 8650, 
    8650, 8650, 8650, 8976, 9375, 9375, 9375, 9375, 9375, 9375,
  8147, 8314, 8095, 8119, 8136, 8149, 8163, 8171, 8180, 8207, 8207, 8207, 
    8207, 8207, 8207, 8767, 9119, 9119, 9119, 9119, 9119, 9119,
  8049, 8223, 7559, 7578, 7591, 7601, 7612, 7619, 7625, 7646, 7646, 7646, 
    7646, 7646, 7646, 8430, 8362, 8362, 8362, 8362, 8362, 8362,
  7742, 7950, 7131, 7155, 7172, 7184, 7198, 7207, 7215, 7241, 7241, 7241, 
    7241, 7241, 7241, 8279, 8138, 8138, 8138, 8138, 8138, 8138,
  6989, 7132, 6361, 6380, 6393, 6404, 6414, 6421, 6429, 6451, 6451, 6451, 
    6451, 6451, 6451, 7881, 7474, 7604, 7604, 7604, 7604, 7604,
  6887, 6900, 5800, 5855, 5894, 5922, 5951, 5969, 5988, 6048, 6048, 6048, 
    6048, 6048, 6048, 7408, 8069, 8069, 8069, 8070, 8069, 8069,
  6658, 6749, 5797, 5843, 5875, 5899, 5923, 5939, 5955, 6006, 6006, 6006, 
    6006, 6006, 6006, 7357, 7706, 7706, 7706, 7706, 7706, 7706,
  6227, 6467, 6263, 6293, 6314, 6330, 6346, 6356, 6368, 6402, 6402, 6402, 
    6402, 6402, 6402, 7570, 7655, 7789, 7789, 7789, 7789, 7789,
  5866, 6139, 6146, 6178, 6201, 6218, 6236, 6247, 6258, 6295, 6295, 6295, 
    6295, 6295, 6295, 7181, 7510, 7510, 7510, 7510, 7510, 7510,
  5642, 5929, 5931, 5968, 5993, 6013, 6033, 6046, 6059, 6099, 6099, 6099, 
    6099, 6099, 6099, 7067, 7473, 7473, 7473, 7473, 7473, 7473,
  5921, 6178, 6023, 6056, 6079, 6096, 6113, 6125, 6137, 6175, 6175, 6175, 
    6175, 6175, 6175, 7374, 7531, 7672, 7672, 7672, 7672, 7672,
  6026, 6230, 5863, 5891, 5911, 5926, 5940, 5950, 5961, 5993, 5993, 5993, 
    5993, 5993, 5993, 7272, 7281, 7424, 7424, 7424, 7424, 7424,
  6132, 6428, 6095, 6137, 6166, 6188, 6211, 6226, 6240, 6287, 6287, 6287, 
    6287, 6287, 6287, 7517, 7853, 7853, 7853, 7853, 7853, 7853,
  5993, 6258, 6010, 6044, 6067, 6085, 6103, 6114, 6127, 6165, 6165, 6165, 
    6165, 6165, 6165, 7485, 7549, 7692, 7692, 7692, 7692, 7692,
  6062, 6297, 5894, 5925, 5947, 5964, 5979, 5990, 6002, 6038, 6038, 6038, 
    6038, 6038, 6038, 7440, 7392, 7537, 7537, 7537, 7537, 7537,
  6314, 6475, 6037, 6097, 6139, 6171, 6202, 6223, 6244, 6311, 6311, 6311, 
    6311, 6311, 6311, 7468, 8543, 8543, 8543, 8543, 8543, 8543,
  6213, 6353, 5938, 5999, 6042, 6073, 6105, 6125, 6147, 6214, 6214, 6214, 
    6214, 6214, 6214, 7280, 8461, 8461, 8461, 8461, 8461, 8461,
  6259, 6410, 6097, 6152, 6190, 6218, 6247, 6265, 6284, 6345, 6345, 6345, 
    6345, 6345, 6345, 7263, 8362, 8362, 8362, 8362, 8362, 8362,
  6354, 6559, 6459, 6498, 6526, 6546, 6567, 6580, 6594, 6637, 6637, 6637, 
    6637, 6637, 6637, 7330, 8093, 8093, 8093, 8093, 8093, 8093,
  6634, 6945, 7141, 7164, 7181, 7193, 7205, 7213, 7221, 7247, 7247, 7247, 
    7247, 7247, 7247, 7778, 8107, 8107, 8107, 8107, 8107, 8107,
  6911, 7230, 7462, 7478, 7489, 7498, 7506, 7511, 7516, 7534, 7534, 7534, 
    7534, 7534, 7534, 7971, 8116, 8116, 8116, 8116, 8116, 8116,
  7281, 7555, 7708, 7718, 7724, 7729, 7734, 7736, 7739, 7749, 7749, 7749, 
    7749, 7749, 7749, 8053, 8082, 8082, 8082, 8082, 8082, 8082,
  7774, 8030, 8167, 8165, 8164, 8163, 8163, 8162, 8161, 8159, 8159, 8159, 
    8159, 8159, 8159, 8311, 8093, 8093, 8093, 8093, 8093, 8093,
  7906, 8142, 8291, 8282, 8275, 8271, 8266, 8262, 8259, 8249, 8249, 8249, 
    8249, 8249, 8249, 8238, 7906, 7906, 7906, 7906, 7906, 7906,
  7773, 8065, 8322, 8313, 8306, 8302, 8297, 8293, 8290, 8280, 8280, 8280, 
    8280, 8280, 8280, 8334, 7935, 7935, 7935, 7935, 7935, 7936,
  7320, 7684, 8097, 8096, 8095, 8094, 8092, 8091, 8091, 8088, 8088, 8088, 
    8088, 8088, 8088, 8276, 8013, 8013, 8013, 8013, 8013, 8013,
  6823, 7180, 7658, 7659, 7660, 7660, 7660, 7660, 7661, 7661, 7661, 7661, 
    7661, 7661, 7661, 7783, 7691, 7691, 7691, 7691, 7691, 7691,
  6349, 6689, 7232, 7233, 7234, 7235, 7236, 7235, 7236, 7237, 7237, 7237, 
    7237, 7237, 7237, 7226, 7271, 7271, 7271, 7271, 7271, 7271,
  6079, 6566, 7412, 7411, 7410, 7410, 7409, 7408, 7408, 7406, 7406, 7406, 
    7406, 7406, 7406, 7509, 7358, 7358, 7357, 7357, 7358, 7358,
  5835, 6431, 7630, 7615, 7606, 7598, 7591, 7585, 7580, 7564, 7564, 7564, 
    7564, 7564, 7564, 7483, 7028, 7028, 7028, 7028, 7028, 7029,
  8776, 8884, 8971, 8974, 8976, 8978, 8980, 8981, 8982, 8986, 8986, 8986, 
    8986, 8986, 8986, 9022, 9106, 9106, 9106, 9106, 9106, 9106,
  8815, 8920, 8992, 8995, 8996, 8998, 9000, 9001, 9002, 9005, 9005, 9005, 
    9005, 9005, 9005, 9034, 9114, 9114, 9114, 9114, 9114, 9114,
  8832, 8936, 9008, 9008, 9007, 9007, 9007, 9007, 9007, 9006, 9006, 9006, 
    9006, 9006, 9006, 9015, 8989, 8989, 8989, 8989, 8989, 8989,
  8843, 8944, 8965, 8967, 8968, 8969, 8971, 8971, 8972, 8974, 8974, 8974, 
    8974, 8974, 8974, 9012, 9044, 9044, 9044, 9044, 9044, 9044,
  8980, 9075, 9100, 9101, 9101, 9101, 9103, 9103, 9103, 9104, 9104, 9104, 
    9104, 9104, 9104, 9110, 9135, 9135, 9135, 9135, 9135, 9135,
  8952, 9045, 9002, 9008, 9012, 9015, 9018, 9020, 9022, 9028, 9028, 9028, 
    9028, 9028, 9028, 9088, 9245, 9245, 9245, 9245, 9245, 9245,
  8957, 9054, 9000, 9005, 9009, 9012, 9016, 9018, 9020, 9026, 9026, 9026, 
    9026, 9026, 9026, 9108, 9245, 9245, 9245, 9245, 9245, 9245,
  8976, 9073, 9051, 9056, 9060, 9062, 9066, 9068, 9070, 9076, 9076, 9076, 
    9076, 9076, 9076, 9139, 9281, 9281, 9281, 9281, 9281, 9281,
  8983, 9080, 9061, 9067, 9072, 9075, 9079, 9081, 9084, 9091, 9091, 9091, 
    9091, 9091, 9091, 9164, 9337, 9337, 9337, 9337, 9337, 9337,
  8956, 9054, 9036, 9044, 9049, 9053, 9058, 9060, 9063, 9071, 9071, 9071, 
    9071, 9071, 9071, 9154, 9356, 9356, 9356, 9356, 9356, 9356,
  8883, 8987, 8852, 8858, 8862, 8864, 8868, 8870, 8872, 8878, 8878, 8878, 
    8878, 8878, 8878, 9034, 9095, 9095, 9095, 9095, 9095, 9095,
  8890, 8990, 8906, 8911, 8915, 8918, 8922, 8923, 8925, 8931, 8931, 8931, 
    8931, 8931, 8931, 9040, 9143, 9143, 9143, 9143, 9143, 9143,
  8911, 9013, 8846, 8851, 8855, 8858, 8861, 8863, 8865, 8871, 8871, 8871, 
    8871, 8871, 8871, 9029, 9072, 9072, 9072, 9072, 9072, 9072,
  9014, 9112, 8984, 8981, 8980, 8979, 8979, 8978, 8977, 8975, 8975, 8975, 
    8975, 8975, 8975, 9053, 8903, 8903, 8903, 8903, 8903, 8903,
  9134, 9222, 9048, 9044, 9040, 9038, 9037, 9035, 9033, 9028, 9028, 9028, 
    9028, 9028, 9028, 9077, 8866, 8866, 8866, 8866, 8866, 8866,
  9218, 9299, 9091, 9082, 9076, 9071, 9068, 9065, 9062, 9052, 9052, 9052, 
    9052, 9052, 9052, 9064, 8738, 8738, 8738, 8738, 8738, 8738,
  9210, 9281, 9005, 8994, 8985, 8979, 8974, 8970, 8966, 8952, 8952, 8952, 
    8952, 8952, 8952, 8940, 8523, 8523, 8523, 8523, 8523, 8523,
  8810, 8918, 8585, 8585, 8585, 8585, 8586, 8586, 8586, 8586, 8586, 8586, 
    8586, 8586, 8586, 8823, 8599, 8599, 8599, 8599, 8599, 8599,
  8971, 9065, 8794, 8790, 8787, 8785, 8784, 8783, 8782, 8777, 8777, 8777, 
    8777, 8777, 8777, 8904, 8642, 8642, 8642, 8642, 8642, 8642,
  8834, 8934, 8688, 8682, 8678, 8675, 8672, 8670, 8668, 8662, 8662, 8662, 
    8662, 8662, 8662, 8787, 8451, 8451, 8451, 8451, 8451, 8451,
  8867, 8968, 8696, 8691, 8688, 8685, 8684, 8682, 8680, 8675, 8675, 8675, 
    8675, 8675, 8675, 8821, 8499, 8499, 8499, 8499, 8499, 8499,
  8886, 8988, 8772, 8769, 8766, 8765, 8764, 8763, 8761, 8757, 8757, 8757, 
    8757, 8757, 8757, 8887, 8638, 8638, 8638, 8638, 8638, 8638,
  8973, 9075, 8799, 8798, 8797, 8796, 8797, 8796, 8796, 8794, 8794, 8794, 
    8794, 8794, 8794, 8976, 8763, 8763, 8763, 8763, 8763, 8763,
  9039, 9135, 8788, 8786, 8784, 8783, 8783, 8783, 8782, 8780, 8780, 8780, 
    8780, 8780, 8780, 8969, 8717, 8717, 8717, 8717, 8717, 8717,
  9193, 9284, 8871, 8869, 8868, 8867, 8866, 8866, 8865, 8862, 8862, 8862, 
    8862, 8862, 8862, 9068, 8790, 8790, 8790, 8790, 8790, 8790,
  9134, 9222, 8809, 8805, 8803, 8801, 8800, 8798, 8797, 8793, 8793, 8793, 
    8793, 8793, 8793, 8971, 8660, 8660, 8660, 8660, 8660, 8660,
  9164, 9252, 8950, 8946, 8943, 8941, 8939, 8938, 8936, 8932, 8932, 8932, 
    8932, 8932, 8932, 9049, 8781, 8781, 8781, 8781, 8781, 8781,
  9300, 9382, 9088, 9083, 9079, 9076, 9074, 9072, 9070, 9063, 9063, 9063, 
    9063, 9063, 9063, 9145, 8860, 8860, 8860, 8860, 8860, 8860,
  9340, 9422, 9057, 9053, 9051, 9049, 9048, 9046, 9045, 9041, 9041, 9041, 
    9041, 9041, 9041, 9172, 8909, 8909, 8909, 8909, 8909, 8909,
  9284, 9369, 8896, 8894, 8893, 8892, 8892, 8891, 8890, 8888, 8888, 8888, 
    8888, 8888, 8888, 9096, 8822, 8822, 8822, 8822, 8822, 8822,
  9232, 9318, 8883, 8881, 8880, 8879, 8879, 8879, 8878, 8876, 8876, 8876, 
    8876, 8876, 8876, 9071, 8824, 8824, 8824, 8824, 8824, 8824,
  9107, 9195, 8835, 8831, 8829, 8827, 8826, 8825, 8824, 8820, 8820, 8820, 
    8820, 8820, 8820, 8971, 8699, 8699, 8699, 8699, 8699, 8699,
  8689, 8804, 8437, 8439, 8441, 8442, 8444, 8445, 8446, 8449, 8449, 8449, 
    8449, 8449, 8449, 8741, 8549, 8549, 8549, 8549, 8549, 8549,
  8345, 8478, 8146, 8151, 8154, 8157, 8161, 8162, 8164, 8170, 8170, 8170, 
    8170, 8170, 8170, 8532, 8367, 8367, 8367, 8367, 8367, 8367,
  8323, 8458, 8064, 8069, 8072, 8075, 8079, 8080, 8082, 8088, 8088, 8088, 
    8088, 8088, 8088, 8488, 8283, 8283, 8283, 8283, 8283, 8283,
  8270, 8405, 8005, 8008, 8011, 8013, 8016, 8018, 8019, 8023, 8023, 8023, 
    8023, 8023, 8023, 8419, 8176, 8176, 8176, 8176, 8176, 8176,
  8359, 8492, 8436, 8442, 8446, 8449, 8453, 8455, 8457, 8464, 8464, 8464, 
    8464, 8464, 8464, 8691, 8695, 8695, 8695, 8695, 8695, 8695,
  8371, 8504, 8452, 8458, 8462, 8465, 8469, 8471, 8473, 8479, 8479, 8479, 
    8479, 8479, 8479, 8699, 8706, 8706, 8706, 8706, 8706, 8706,
  8376, 8503, 8278, 8281, 8283, 8285, 8288, 8289, 8290, 8293, 8293, 8293, 
    8293, 8293, 8293, 8564, 8423, 8423, 8423, 8423, 8423, 8423,
  8366, 8491, 8260, 8262, 8263, 8264, 8266, 8267, 8268, 8270, 8270, 8270, 
    8270, 8270, 8270, 8527, 8358, 8358, 8358, 8358, 8358, 8358,
  8263, 8395, 8217, 8220, 8223, 8225, 8228, 8229, 8230, 8234, 8234, 8234, 
    8234, 8234, 8234, 8499, 8379, 8379, 8379, 8379, 8379, 8379,
  8000, 8144, 8026, 8030, 8033, 8035, 8038, 8040, 8041, 8046, 8046, 8046, 
    8046, 8046, 8046, 8331, 8213, 8213, 8213, 8213, 8213, 8213,
  8073, 8221, 8233, 8242, 8248, 8253, 8258, 8262, 8265, 8275, 8275, 8275, 
    8275, 8275, 8275, 8543, 8621, 8621, 8621, 8621, 8621, 8621,
  8015, 8167, 8120, 8131, 8138, 8144, 8150, 8154, 8158, 8170, 8170, 8170, 
    8170, 8170, 8170, 8490, 8577, 8577, 8577, 8577, 8577, 8577,
  7965, 8118, 8098, 8108, 8115, 8120, 8127, 8130, 8134, 8145, 8145, 8145, 
    8145, 8145, 8145, 8454, 8530, 8530, 8530, 8530, 8530, 8530,
  7897, 8054, 8118, 8128, 8135, 8140, 8146, 8149, 8153, 8163, 8163, 8163, 
    8163, 8163, 8163, 8441, 8535, 8535, 8535, 8535, 8535, 8535,
  8007, 8157, 8159, 8168, 8175, 8180, 8186, 8189, 8192, 8202, 8202, 8202, 
    8202, 8202, 8202, 8480, 8555, 8555, 8555, 8555, 8555, 8555,
  8177, 8316, 8216, 8224, 8229, 8233, 8238, 8240, 8243, 8251, 8251, 8251, 
    8251, 8251, 8251, 8529, 8539, 8539, 8539, 8539, 8539, 8539,
  8325, 8455, 8327, 8333, 8336, 8339, 8343, 8345, 8347, 8352, 8352, 8352, 
    8352, 8352, 8352, 8599, 8560, 8560, 8560, 8560, 8560, 8560,
  8386, 8513, 8383, 8388, 8391, 8394, 8397, 8399, 8401, 8406, 8406, 8406, 
    8406, 8406, 8406, 8640, 8604, 8604, 8604, 8604, 8604, 8604,
  8345, 8475, 8351, 8356, 8360, 8362, 8366, 8368, 8370, 8375, 8375, 8375, 
    8375, 8375, 8375, 8616, 8577, 8577, 8577, 8577, 8577, 8577,
  8144, 8271, 7954, 7955, 7956, 7957, 7958, 7959, 7959, 7960, 7960, 7960, 
    7960, 7960, 7960, 8255, 8016, 8016, 8016, 8016, 8016, 8016,
  8108, 8241, 8029, 8030, 8030, 8031, 8033, 8033, 8033, 8034, 8034, 8034, 
    8034, 8034, 8034, 8303, 8081, 8081, 8081, 8081, 8081, 8081,
  8043, 8192, 7897, 7900, 7902, 7903, 7906, 7907, 7908, 7910, 7910, 7910, 
    7910, 7910, 7910, 8298, 8021, 8021, 8021, 8021, 8021, 8021,
  7924, 8088, 7733, 7745, 7754, 7761, 7768, 7773, 7777, 7791, 7791, 7791, 
    7791, 7791, 7791, 8334, 8271, 8271, 8271, 8271, 8271, 8271,
  7748, 7919, 7535, 7547, 7555, 7561, 7568, 7573, 7577, 7590, 7590, 7590, 
    7590, 7590, 7590, 8166, 8040, 8040, 8040, 8040, 8040, 8040,
  7586, 7767, 7334, 7353, 7366, 7376, 7387, 7394, 7400, 7422, 7422, 7422, 
    7422, 7422, 7422, 8103, 8142, 8142, 8142, 8142, 8142, 8142,
  7445, 7633, 7212, 7234, 7249, 7261, 7273, 7281, 7289, 7313, 7313, 7313, 
    7313, 7313, 7313, 8032, 8134, 8134, 8134, 8134, 8134, 8134,
  7433, 7627, 7271, 7290, 7303, 7313, 7324, 7331, 7337, 7359, 7359, 7359, 
    7359, 7359, 7359, 8055, 8076, 8076, 8076, 8076, 8076, 8076,
  7490, 7679, 7376, 7393, 7405, 7415, 7425, 7431, 7437, 7457, 7457, 7457, 
    7457, 7457, 7457, 8099, 8120, 8120, 8120, 8120, 8120, 8120,
  7619, 7809, 7556, 7570, 7580, 7587, 7596, 7601, 7605, 7621, 7621, 7621, 
    7621, 7621, 7621, 8226, 8149, 8149, 8149, 8149, 8149, 8149,
  7658, 7841, 7771, 7785, 7794, 7801, 7809, 7814, 7819, 7834, 7834, 7834, 
    7834, 7834, 7834, 8311, 8344, 8344, 8344, 8344, 8344, 8344,
  7735, 7924, 8121, 8141, 8155, 8165, 8177, 8184, 8191, 8213, 8213, 8213, 
    8213, 8213, 8213, 8622, 8969, 8969, 8968, 8968, 8968, 8969,
  7765, 7948, 8195, 8216, 8231, 8242, 8254, 8262, 8269, 8293, 8293, 8293, 
    8293, 8293, 8293, 8655, 9099, 9099, 9099, 9099, 9099, 9099,
  7826, 8012, 8186, 8211, 8229, 8243, 8258, 8266, 8276, 8304, 8304, 8304, 
    8304, 8304, 8304, 8747, 9274, 9274, 9274, 9274, 9274, 9274,
  7785, 7982, 7992, 8025, 8047, 8064, 8082, 8093, 8105, 8141, 8141, 8141, 
    8141, 8141, 8141, 8756, 9356, 9356, 9356, 9356, 9356, 9356,
  7729, 7922, 7584, 7620, 7646, 7665, 7685, 7698, 7711, 7752, 7752, 7752, 
    7752, 7752, 7752, 8550, 9125, 9125, 9125, 9125, 9125, 9125,
  7871, 8048, 7362, 7382, 7396, 7407, 7418, 7426, 7433, 7455, 7455, 7455, 
    7455, 7455, 7455, 8271, 8220, 8220, 8220, 8220, 8220, 8220,
  7394, 7526, 7043, 7058, 7069, 7077, 7086, 7091, 7097, 7115, 7115, 7115, 
    7115, 7115, 7115, 8131, 7914, 8023, 8023, 8023, 8023, 8023,
  6970, 7125, 6679, 6699, 6712, 6723, 6733, 6740, 6748, 6770, 6770, 6770, 
    6770, 6770, 6770, 7871, 7727, 7848, 7848, 7848, 7848, 7848,
  6859, 6978, 6289, 6336, 6369, 6393, 6417, 6433, 6450, 6501, 6501, 6501, 
    6501, 6501, 6501, 7655, 8224, 8224, 8224, 8224, 8224, 8224,
  6496, 6622, 5887, 5936, 5970, 5995, 6020, 6036, 6053, 6106, 6106, 6106, 
    6106, 6106, 6106, 7353, 7891, 7890, 7891, 7891, 7890, 7891,
  6221, 6336, 5521, 5579, 5619, 5649, 5679, 5699, 5719, 5783, 5783, 5783, 
    5783, 5783, 5783, 7183, 7916, 7915, 7915, 7916, 7915, 7915,
  5830, 6056, 5679, 5710, 5732, 5749, 5765, 5775, 5787, 5823, 5823, 5823, 
    5823, 5823, 5823, 7204, 7216, 7366, 7366, 7366, 7366, 7366,
  5656, 5912, 5705, 5739, 5763, 5782, 5799, 5811, 5824, 5863, 5863, 5863, 
    5863, 5863, 5863, 7158, 7308, 7457, 7457, 7457, 7457, 7457,
  5559, 5814, 5627, 5661, 5685, 5703, 5721, 5733, 5746, 5786, 5786, 5786, 
    5786, 5786, 5786, 7070, 7248, 7400, 7400, 7400, 7400, 7400,
  5633, 5904, 5623, 5659, 5684, 5703, 5722, 5734, 5748, 5789, 5789, 5789, 
    5789, 5789, 5789, 7213, 7296, 7450, 7450, 7450, 7450, 7450,
  5577, 5801, 5396, 5428, 5451, 5468, 5484, 5496, 5508, 5545, 5545, 5545, 
    5545, 5545, 5545, 6985, 7009, 7167, 7167, 7167, 7167, 7167,
  5569, 5831, 5486, 5521, 5546, 5566, 5584, 5596, 5610, 5651, 5651, 5651, 
    5651, 5651, 5651, 7134, 7178, 7335, 7335, 7335, 7335, 7335,
  5564, 5833, 5565, 5601, 5626, 5646, 5664, 5676, 5690, 5731, 5731, 5731, 
    5731, 5731, 5731, 7142, 7247, 7402, 7402, 7402, 7402, 7402,
  5517, 5762, 5440, 5474, 5498, 5516, 5534, 5546, 5559, 5598, 5598, 5598, 
    5598, 5598, 5598, 7015, 7099, 7257, 7257, 7257, 7257, 7257,
  5553, 5789, 5455, 5487, 5511, 5529, 5546, 5557, 5570, 5608, 5608, 5608, 
    5608, 5608, 5608, 7006, 7084, 7241, 7241, 7241, 7241, 7241,
  5620, 5843, 5795, 5825, 5847, 5863, 5879, 5890, 5902, 5937, 5937, 5937, 
    5937, 5937, 5937, 6969, 7278, 7421, 7421, 7421, 7421, 7421,
  6139, 6362, 6266, 6312, 6344, 6368, 6391, 6407, 6423, 6473, 6473, 6473, 
    6473, 6473, 6473, 7287, 8164, 8164, 8164, 8164, 8164, 8164,
  6369, 6603, 6982, 7008, 7027, 7042, 7056, 7065, 7075, 7105, 7105, 7105, 
    7105, 7105, 7105, 7576, 8126, 8236, 8236, 8236, 8236, 8236,
  6730, 6978, 7426, 7452, 7471, 7485, 7499, 7508, 7518, 7547, 7547, 7547, 
    7547, 7547, 7547, 7926, 8474, 8573, 8573, 8573, 8573, 8573,
  7080, 7410, 7679, 7692, 7701, 7708, 7714, 7718, 7723, 7737, 7737, 7737, 
    7737, 7737, 7737, 8135, 8209, 8209, 8209, 8209, 8209, 8209,
  7442, 7678, 7759, 7768, 7775, 7779, 7784, 7786, 7790, 7799, 7799, 7799, 
    7799, 7799, 7799, 8062, 8124, 8124, 8124, 8124, 8124, 8124,
  7903, 8112, 8143, 8142, 8141, 8140, 8140, 8139, 8138, 8137, 8137, 8137, 
    8137, 8137, 8137, 8257, 8082, 8081, 8081, 8082, 8082, 8082,
  8052, 8244, 8281, 8274, 8269, 8265, 8261, 8258, 8255, 8247, 8247, 8247, 
    8247, 8247, 8247, 8243, 7969, 7969, 7969, 7969, 7969, 7969,
  7913, 8168, 8362, 8354, 8349, 8345, 8341, 8338, 8335, 8326, 8326, 8326, 
    8326, 8326, 8326, 8344, 8036, 8036, 8036, 8036, 8036, 8036,
  7446, 7787, 8182, 8177, 8174, 8171, 8168, 8166, 8164, 8158, 8158, 8158, 
    8158, 8158, 8158, 8256, 7961, 7961, 7961, 7961, 7961, 7961,
  6944, 7284, 7726, 7726, 7726, 7726, 7726, 7725, 7725, 7725, 7725, 7725, 
    7725, 7725, 7725, 7821, 7720, 7720, 7720, 7720, 7720, 7720,
  6540, 6842, 7275, 7277, 7279, 7281, 7282, 7282, 7283, 7285, 7285, 7285, 
    7285, 7285, 7285, 7291, 7368, 7368, 7368, 7368, 7368, 7368,
  6145, 6574, 7317, 7317, 7317, 7316, 7316, 7315, 7315, 7315, 7315, 7315, 
    7315, 7315, 7315, 7356, 7295, 7295, 7295, 7295, 7296, 7296,
  6059, 6598, 7560, 7556, 7553, 7551, 7548, 7546, 7545, 7539, 7539, 7539, 
    7539, 7539, 7539, 7646, 7368, 7368, 7368, 7368, 7369, 7369,
  8745, 8853, 8981, 8984, 8987, 8989, 8992, 8993, 8994, 8998, 8998, 8998, 
    8998, 8998, 8998, 9019, 9144, 9144, 9144, 9144, 9144, 9144,
  8791, 8897, 8955, 8957, 8958, 8959, 8961, 8962, 8962, 8964, 8964, 8964, 
    8964, 8964, 8964, 8999, 9040, 9040, 9040, 9040, 9040, 9040,
  8813, 8917, 8971, 8973, 8975, 8976, 8978, 8979, 8980, 8982, 8982, 8982, 
    8982, 8982, 8982, 9015, 9071, 9071, 9071, 9071, 9071, 9071,
  8865, 8969, 9033, 9033, 9034, 9034, 9035, 9036, 9036, 9037, 9037, 9037, 
    9037, 9037, 9037, 9057, 9072, 9072, 9072, 9072, 9072, 9072,
  8945, 9042, 9040, 9042, 9044, 9045, 9047, 9048, 9049, 9051, 9051, 9051, 
    9051, 9051, 9051, 9090, 9147, 9147, 9147, 9147, 9147, 9147,
  8999, 9090, 9147, 9151, 9153, 9155, 9157, 9158, 9160, 9163, 9163, 9163, 
    9163, 9163, 9163, 9153, 9298, 9298, 9297, 9297, 9298, 9298,
  8922, 9015, 8974, 8980, 8984, 8987, 8990, 8992, 8994, 9000, 9000, 9000, 
    9000, 9000, 9000, 9059, 9215, 9215, 9215, 9215, 9215, 9215,
  8917, 9018, 8986, 8991, 8994, 8997, 9000, 9002, 9004, 9009, 9009, 9009, 
    9009, 9009, 9009, 9092, 9205, 9205, 9205, 9205, 9205, 9205,
  8934, 9034, 8991, 8996, 9000, 9003, 9006, 9008, 9010, 9016, 9016, 9016, 
    9016, 9016, 9016, 9107, 9221, 9221, 9221, 9221, 9221, 9221,
  8998, 9100, 9043, 9048, 9051, 9053, 9056, 9058, 9060, 9065, 9065, 9065, 
    9065, 9065, 9065, 9168, 9243, 9243, 9243, 9243, 9243, 9243,
  8971, 9073, 9003, 9006, 9008, 9009, 9012, 9013, 9014, 9017, 9017, 9017, 
    9017, 9017, 9017, 9114, 9134, 9134, 9134, 9134, 9134, 9134,
  9040, 9140, 9051, 9049, 9048, 9047, 9047, 9046, 9046, 9044, 9044, 9044, 
    9044, 9044, 9044, 9120, 8992, 8992, 8992, 8992, 8992, 8992,
  8989, 9091, 8970, 8970, 8969, 8969, 8970, 8970, 8970, 8969, 8969, 8969, 
    8969, 8969, 8969, 9073, 8967, 8967, 8967, 8967, 8967, 8967,
  9016, 9110, 8940, 8937, 8936, 8934, 8934, 8933, 8932, 8929, 8929, 8929, 
    8929, 8929, 8929, 9011, 8843, 8843, 8843, 8843, 8843, 8843,
  9140, 9218, 8936, 8927, 8921, 8916, 8913, 8910, 8907, 8897, 8897, 8897, 
    8897, 8897, 8897, 8938, 8586, 8586, 8586, 8586, 8586, 8586,
  9089, 9168, 8848, 8838, 8831, 8826, 8822, 8818, 8814, 8803, 8803, 8803, 
    8803, 8803, 8803, 8855, 8439, 8439, 8439, 8439, 8439, 8439,
  9014, 9106, 8831, 8826, 8823, 8820, 8819, 8817, 8815, 8810, 8810, 8810, 
    8810, 8810, 8810, 8924, 8643, 8643, 8643, 8643, 8643, 8643,
  9010, 9101, 8804, 8800, 8797, 8795, 8794, 8792, 8791, 8786, 8786, 8786, 
    8786, 8786, 8786, 8912, 8640, 8640, 8640, 8640, 8640, 8640,
  8990, 9084, 8884, 8879, 8876, 8874, 8873, 8871, 8870, 8865, 8865, 8865, 
    8865, 8865, 8865, 8953, 8713, 8713, 8713, 8713, 8713, 8713,
  8983, 9082, 8803, 8801, 8800, 8799, 8799, 8798, 8797, 8795, 8795, 8795, 
    8795, 8795, 8795, 8960, 8735, 8735, 8735, 8735, 8735, 8735,
  9044, 9137, 8832, 8827, 8823, 8820, 8817, 8815, 8813, 8807, 8807, 8807, 
    8807, 8807, 8807, 8937, 8601, 8601, 8601, 8601, 8601, 8601,
  8912, 9016, 8788, 8786, 8785, 8784, 8784, 8783, 8782, 8780, 8780, 8780, 
    8780, 8780, 8780, 8938, 8720, 8720, 8720, 8720, 8720, 8720,
  8873, 8978, 8827, 8828, 8828, 8828, 8830, 8830, 8830, 8830, 8830, 8830, 
    8830, 8830, 8830, 8964, 8859, 8859, 8859, 8859, 8859, 8859,
  9033, 9134, 8699, 8699, 8698, 8698, 8699, 8699, 8699, 8699, 8699, 8699, 
    8699, 8699, 8699, 8968, 8708, 8708, 8708, 8708, 8708, 8708,
  9131, 9221, 8791, 8788, 8786, 8785, 8784, 8783, 8782, 8779, 8779, 8779, 
    8779, 8779, 8779, 8980, 8681, 8681, 8681, 8681, 8681, 8681,
  9229, 9315, 9018, 9014, 9012, 9009, 9008, 9007, 9006, 9001, 9001, 9001, 
    9001, 9001, 9001, 9114, 8862, 8862, 8862, 8862, 8862, 8862,
  9167, 9257, 8882, 8880, 8879, 8878, 8878, 8877, 8876, 8874, 8874, 8874, 
    8874, 8874, 8874, 9052, 8809, 8809, 8809, 8809, 8809, 8809,
  9301, 9383, 9030, 9027, 9025, 9023, 9022, 9021, 9020, 9017, 9017, 9017, 
    9017, 9017, 9017, 9152, 8913, 8913, 8913, 8913, 8913, 8913,
  9383, 9461, 9049, 9045, 9042, 9040, 9039, 9037, 9036, 9031, 9031, 9031, 
    9031, 9031, 9031, 9172, 8891, 8891, 8891, 8891, 8891, 8891,
  9313, 9393, 8943, 8940, 8938, 8936, 8935, 8934, 8932, 8929, 8929, 8929, 
    8929, 8929, 8929, 9101, 8810, 8810, 8810, 8810, 8810, 8810,
  9293, 9372, 8952, 8948, 8946, 8944, 8943, 8942, 8940, 8936, 8936, 8936, 
    8936, 8936, 8936, 9088, 8813, 8813, 8813, 8813, 8813, 8813,
  9265, 9348, 8946, 8944, 8942, 8941, 8941, 8940, 8939, 8937, 8937, 8937, 
    8937, 8937, 8937, 9096, 8859, 8859, 8859, 8859, 8859, 8859,
  8988, 9084, 8725, 8724, 8723, 8722, 8723, 8722, 8722, 8720, 8720, 8720, 
    8720, 8720, 8720, 8916, 8682, 8682, 8682, 8682, 8682, 8682,
  8931, 9030, 8710, 8710, 8710, 8710, 8710, 8710, 8710, 8710, 8710, 8710, 
    8710, 8710, 8710, 8903, 8706, 8706, 8706, 8706, 8706, 8706,
  8423, 8551, 8188, 8192, 8194, 8196, 8199, 8200, 8202, 8206, 8206, 8206, 
    8206, 8206, 8206, 8552, 8350, 8350, 8350, 8350, 8350, 8350,
  8447, 8576, 8229, 8234, 8237, 8240, 8243, 8245, 8246, 8252, 8252, 8252, 
    8252, 8252, 8252, 8604, 8435, 8435, 8435, 8435, 8435, 8435,
  8400, 8530, 8120, 8125, 8129, 8132, 8135, 8137, 8139, 8144, 8144, 8144, 
    8144, 8144, 8144, 8533, 8341, 8341, 8341, 8341, 8341, 8341,
  8236, 8370, 8078, 8081, 8083, 8084, 8087, 8088, 8089, 8092, 8092, 8092, 
    8092, 8092, 8092, 8420, 8212, 8212, 8212, 8212, 8212, 8212,
  8336, 8467, 8210, 8214, 8217, 8219, 8222, 8224, 8225, 8229, 8229, 8229, 
    8229, 8229, 8229, 8538, 8394, 8394, 8394, 8394, 8394, 8394,
  8237, 8375, 8228, 8232, 8235, 8238, 8241, 8242, 8244, 8249, 8249, 8249, 
    8249, 8249, 8249, 8533, 8424, 8424, 8424, 8424, 8424, 8424,
  8326, 8457, 8220, 8223, 8225, 8227, 8230, 8231, 8232, 8235, 8235, 8235, 
    8235, 8235, 8235, 8523, 8361, 8361, 8361, 8361, 8361, 8361,
  8126, 8262, 8026, 8029, 8031, 8033, 8035, 8036, 8037, 8040, 8040, 8040, 
    8040, 8040, 8040, 8342, 8162, 8162, 8162, 8162, 8162, 8162,
  7985, 8127, 7956, 7960, 7963, 7965, 7969, 7970, 7971, 7976, 7976, 7976, 
    7976, 7976, 7976, 8274, 8138, 8138, 8138, 8138, 8138, 8138,
  7994, 8145, 8134, 8143, 8150, 8155, 8161, 8164, 8167, 8178, 8178, 8178, 
    8178, 8178, 8178, 8469, 8539, 8539, 8539, 8539, 8539, 8539,
  8003, 8154, 8070, 8080, 8087, 8092, 8098, 8102, 8105, 8116, 8116, 8116, 
    8116, 8116, 8116, 8448, 8490, 8490, 8490, 8490, 8490, 8490,
  7927, 8082, 8095, 8105, 8111, 8117, 8123, 8126, 8129, 8140, 8140, 8140, 
    8140, 8140, 8140, 8433, 8510, 8510, 8510, 8510, 8510, 8510,
  7985, 8136, 8161, 8170, 8177, 8181, 8187, 8190, 8193, 8204, 8204, 8204, 
    8204, 8204, 8204, 8473, 8551, 8551, 8551, 8551, 8551, 8551,
  8218, 8355, 8258, 8264, 8269, 8272, 8276, 8278, 8280, 8287, 8287, 8287, 
    8287, 8287, 8287, 8547, 8524, 8524, 8524, 8524, 8524, 8524,
  8331, 8462, 8311, 8316, 8320, 8323, 8327, 8329, 8330, 8336, 8336, 8336, 
    8336, 8336, 8336, 8595, 8543, 8543, 8543, 8543, 8543, 8543,
  8409, 8535, 8368, 8373, 8376, 8379, 8382, 8384, 8386, 8391, 8391, 8391, 
    8391, 8391, 8391, 8639, 8581, 8581, 8581, 8581, 8581, 8581,
  8380, 8507, 8361, 8366, 8369, 8372, 8375, 8377, 8379, 8384, 8384, 8384, 
    8384, 8384, 8384, 8624, 8570, 8570, 8570, 8570, 8570, 8570,
  8367, 8489, 8195, 8196, 8196, 8196, 8197, 8197, 8197, 8197, 8197, 8197, 
    8197, 8197, 8197, 8458, 8211, 8211, 8211, 8211, 8211, 8211,
  8127, 8266, 7948, 7951, 7952, 7953, 7956, 7957, 7957, 7960, 7960, 7960, 
    7960, 7960, 7960, 8316, 8054, 8054, 8054, 8054, 8054, 8054,
  8141, 8283, 8117, 8123, 8127, 8130, 8134, 8136, 8138, 8145, 8145, 8145, 
    8145, 8145, 8145, 8460, 8380, 8380, 8380, 8380, 8380, 8380,
  8127, 8282, 7657, 7670, 7679, 7686, 7694, 7699, 7704, 7718, 7718, 7718, 
    7718, 7718, 7718, 8367, 8218, 8218, 8218, 8218, 8218, 8218,
  7900, 8060, 7510, 7524, 7534, 7542, 7550, 7555, 7560, 7576, 7576, 7576, 
    7576, 7576, 7576, 8209, 8122, 8122, 8122, 8122, 8122, 8122,
  7550, 7729, 7376, 7395, 7408, 7418, 7429, 7436, 7443, 7464, 7464, 7464, 
    7464, 7464, 7464, 8095, 8178, 8178, 8178, 8178, 8178, 8178,
  7364, 7561, 7194, 7214, 7229, 7240, 7252, 7259, 7267, 7290, 7290, 7290, 
    7290, 7290, 7290, 8014, 8075, 8075, 8075, 8075, 8075, 8075,
  7239, 7448, 7084, 7104, 7118, 7129, 7141, 7148, 7155, 7177, 7177, 7177, 
    7177, 7177, 7177, 7947, 7943, 7943, 7943, 7943, 7943, 7943,
  6989, 7205, 6937, 6960, 6976, 6988, 7001, 7009, 7017, 7042, 7042, 7042, 
    7042, 7042, 7042, 7802, 7899, 7899, 7899, 7899, 7899, 7899,
  6950, 7177, 6862, 6884, 6899, 6911, 6924, 6932, 6939, 6964, 6964, 6964, 
    6964, 6964, 6964, 7790, 7804, 7804, 7804, 7804, 7804, 7804,
  6960, 7190, 6755, 6779, 6795, 6808, 6822, 6830, 6838, 6865, 6865, 6865, 
    6865, 6865, 6865, 7776, 7765, 7765, 7765, 7765, 7765, 7765,
  6849, 7075, 7048, 7073, 7091, 7105, 7118, 7126, 7137, 7165, 7165, 7165, 
    7165, 7165, 7165, 8005, 8162, 8273, 8273, 8273, 8273, 8273,
  7075, 7296, 6759, 6785, 6803, 6817, 6832, 6841, 6850, 6879, 6879, 6879, 
    6879, 6879, 6879, 7822, 7867, 7867, 7867, 7867, 7867, 7867,
  7264, 7486, 6831, 6857, 6874, 6888, 6902, 6911, 6920, 6948, 6948, 6948, 
    6948, 6948, 6948, 7958, 7901, 7901, 7901, 7901, 7901, 7901,
  7062, 7273, 6968, 6991, 7008, 7021, 7033, 7041, 7051, 7078, 7078, 7078, 
    7078, 7078, 7078, 8158, 8074, 8189, 8189, 8189, 8189, 8189,
  7131, 7308, 6879, 6899, 6914, 6925, 6936, 6943, 6951, 6975, 6975, 6975, 
    6975, 6975, 6975, 8094, 7923, 8039, 8039, 8039, 8039, 8039,
  7053, 7213, 6796, 6815, 6829, 6839, 6849, 6856, 6864, 6886, 6886, 6886, 
    6886, 6886, 6886, 7955, 7817, 7934, 7934, 7934, 7934, 7934,
  6944, 7111, 6791, 6811, 6825, 6836, 6847, 6854, 6862, 6885, 6885, 6885, 
    6885, 6885, 6885, 7881, 7834, 7952, 7952, 7952, 7952, 7952,
  6675, 6888, 6753, 6778, 6796, 6809, 6822, 6831, 6841, 6869, 6869, 6869, 
    6869, 6869, 6869, 7820, 7923, 8042, 8042, 8042, 8042, 8042,
  6329, 6548, 6416, 6444, 6463, 6478, 6492, 6501, 6512, 6543, 6543, 6543, 
    6543, 6543, 6543, 7559, 7710, 7839, 7839, 7839, 7839, 7839,
  6066, 6300, 6160, 6189, 6210, 6227, 6242, 6252, 6264, 6298, 6298, 6298, 
    6298, 6298, 6298, 7401, 7567, 7703, 7703, 7703, 7703, 7703,
  5782, 5995, 5715, 5744, 5765, 5782, 5797, 5807, 5819, 5853, 5853, 5853, 
    5853, 5853, 5853, 7096, 7203, 7351, 7351, 7351, 7351, 7351,
  5650, 5868, 5470, 5501, 5523, 5540, 5556, 5567, 5579, 5615, 5615, 5615, 
    5615, 5615, 5615, 7021, 7047, 7202, 7202, 7202, 7202, 7202,
  5594, 5842, 5464, 5498, 5522, 5541, 5558, 5570, 5583, 5623, 5623, 5623, 
    5623, 5623, 5623, 7098, 7123, 7279, 7279, 7279, 7279, 7279,
  5502, 5763, 5451, 5486, 5511, 5530, 5548, 5561, 5574, 5615, 5615, 5615, 
    5615, 5615, 5615, 7068, 7148, 7306, 7306, 7306, 7306, 7306,
  5307, 5552, 5167, 5201, 5226, 5245, 5263, 5276, 5289, 5330, 5330, 5330, 
    5330, 5330, 5330, 6844, 6906, 7070, 7070, 7070, 7070, 7070,
  5209, 5462, 5202, 5237, 5263, 5282, 5301, 5313, 5327, 5368, 5368, 5368, 
    5368, 5368, 5368, 6780, 6950, 7113, 7113, 7113, 7113, 7113,
  5155, 5428, 5268, 5305, 5332, 5352, 5372, 5385, 5399, 5443, 5443, 5443, 
    5443, 5443, 5443, 6802, 7048, 7210, 7210, 7210, 7210, 7210,
  5123, 5395, 5255, 5293, 5319, 5339, 5359, 5372, 5386, 5430, 5430, 5430, 
    5430, 5430, 5430, 6771, 7035, 7197, 7197, 7197, 7197, 7197,
  5154, 5432, 5286, 5324, 5351, 5371, 5391, 5404, 5419, 5463, 5463, 5463, 
    5463, 5463, 5463, 6825, 7078, 7240, 7240, 7240, 7240, 7240,
  5319, 5580, 5407, 5442, 5468, 5487, 5506, 5518, 5532, 5573, 5573, 5573, 
    5573, 5573, 5573, 6895, 7117, 7275, 7275, 7275, 7275, 7275,
  5667, 5908, 5719, 5751, 5774, 5792, 5809, 5820, 5833, 5870, 5870, 5870, 
    5870, 5870, 5870, 7103, 7279, 7428, 7428, 7428, 7428, 7428,
  6107, 6338, 6571, 6599, 6619, 6634, 6649, 6658, 6670, 6702, 6702, 6702, 
    6702, 6702, 6702, 7368, 7835, 7957, 7957, 7957, 7957, 7957,
  6632, 6892, 7344, 7372, 7392, 7407, 7421, 7431, 7442, 7473, 7473, 7473, 
    7473, 7473, 7473, 7895, 8451, 8552, 8552, 8552, 8552, 8552,
  7037, 7393, 7712, 7725, 7734, 7741, 7748, 7752, 7757, 7771, 7771, 7771, 
    7771, 7771, 7771, 8205, 8256, 8256, 8256, 8256, 8256, 8256,
  7385, 7694, 7840, 7851, 7859, 7865, 7871, 7874, 7878, 7890, 7890, 7890, 
    7890, 7890, 7890, 8340, 8295, 8295, 8295, 8295, 8295, 8295,
  7718, 7925, 7868, 7878, 7886, 7891, 7897, 7900, 7903, 7915, 7915, 7915, 
    7915, 7915, 7915, 8255, 8299, 8299, 8299, 8299, 8299, 8299,
  8079, 8157, 8184, 8182, 8182, 8180, 8179, 8178, 8179, 8176, 8176, 8176, 
    8176, 8176, 8176, 8098, 8107, 8107, 8107, 8107, 8107, 8107,
  8084, 8237, 8388, 8377, 8371, 8365, 8359, 8355, 8353, 8340, 8340, 8340, 
    8340, 8340, 8340, 8190, 7953, 7953, 7953, 7953, 7953, 7953,
  7978, 8257, 8495, 8484, 8477, 8471, 8465, 8461, 8457, 8445, 8445, 8445, 
    8445, 8445, 8445, 8457, 8036, 8036, 8036, 8036, 8036, 8036,
  7578, 7912, 8291, 8283, 8278, 8274, 8270, 8267, 8264, 8255, 8255, 8255, 
    8255, 8255, 8255, 8323, 7966, 7966, 7966, 7966, 7966, 7966,
  7144, 7496, 7962, 7957, 7955, 7952, 7950, 7948, 7946, 7941, 7941, 7941, 
    7941, 7941, 7941, 7998, 7770, 7770, 7770, 7770, 7770, 7770,
  6730, 7026, 7465, 7464, 7463, 7463, 7462, 7461, 7461, 7459, 7459, 7459, 
    7459, 7459, 7459, 7402, 7414, 7414, 7413, 7413, 7414, 7414,
  6410, 6802, 7452, 7450, 7448, 7447, 7445, 7444, 7443, 7439, 7439, 7439, 
    7439, 7439, 7439, 7436, 7330, 7330, 7330, 7330, 7330, 7330,
  6184, 6698, 7613, 7606, 7601, 7598, 7594, 7591, 7588, 7580, 7580, 7580, 
    7580, 7580, 7580, 7630, 7315, 7315, 7315, 7315, 7315, 7316,
  8725, 8832, 8963, 8964, 8964, 8965, 8966, 8967, 8967, 8968, 8968, 8968, 
    8968, 8968, 8968, 8965, 9019, 9019, 9019, 9019, 9019, 9019,
  8823, 8929, 9028, 9028, 9028, 9028, 9029, 9029, 9029, 9029, 9029, 9029, 
    9029, 9029, 9029, 9034, 9048, 9048, 9048, 9048, 9048, 9048,
  8817, 8921, 8975, 8977, 8978, 8978, 8980, 8980, 8981, 8982, 8982, 8982, 
    8982, 8982, 8982, 9010, 9038, 9038, 9038, 9038, 9038, 9038,
  8896, 8999, 9034, 9035, 9037, 9038, 9040, 9040, 9041, 9043, 9043, 9043, 
    9043, 9043, 9043, 9086, 9124, 9124, 9124, 9124, 9124, 9124,
  8975, 9073, 9105, 9104, 9104, 9104, 9104, 9104, 9104, 9103, 9103, 9103, 
    9103, 9103, 9103, 9114, 9095, 9095, 9095, 9095, 9095, 9095,
  9022, 9112, 9152, 9156, 9158, 9160, 9163, 9164, 9165, 9169, 9169, 9169, 
    9169, 9169, 9169, 9162, 9310, 9310, 9310, 9310, 9310, 9310,
  8943, 9039, 9001, 9005, 9008, 9010, 9013, 9014, 9016, 9020, 9020, 9020, 
    9020, 9020, 9020, 9082, 9182, 9182, 9182, 9182, 9182, 9182,
  8916, 9013, 9016, 9020, 9024, 9026, 9029, 9031, 9032, 9037, 9037, 9037, 
    9037, 9037, 9037, 9082, 9214, 9214, 9214, 9214, 9214, 9214,
  8852, 8954, 8907, 8911, 8914, 8916, 8920, 8921, 8923, 8927, 8927, 8927, 
    8927, 8927, 8927, 9020, 9099, 9099, 9099, 9099, 9099, 9099,
  8935, 9037, 8989, 8990, 8992, 8992, 8994, 8995, 8995, 8997, 8997, 8997, 
    8997, 8997, 8997, 9076, 9067, 9067, 9067, 9067, 9067, 9067,
  8990, 9092, 8999, 8998, 8998, 8997, 8997, 8997, 8997, 8996, 8996, 8996, 
    8996, 8996, 8996, 9084, 8967, 8967, 8967, 8967, 8967, 8967,
  8964, 9066, 8972, 8972, 8971, 8971, 8971, 8971, 8971, 8970, 8970, 8970, 
    8970, 8970, 8970, 9059, 8952, 8952, 8952, 8952, 8952, 8952,
  9008, 9104, 8971, 8969, 8967, 8965, 8965, 8964, 8963, 8960, 8960, 8960, 
    8960, 8960, 8960, 9028, 8867, 8867, 8867, 8867, 8867, 8867,
  9222, 9296, 9087, 9077, 9070, 9065, 9060, 9057, 9053, 9042, 9042, 9042, 
    9042, 9042, 9042, 9024, 8683, 8683, 8683, 8683, 8683, 8683,
  8956, 9046, 8768, 8763, 8760, 8757, 8756, 8754, 8752, 8747, 8747, 8747, 
    8747, 8747, 8747, 8852, 8577, 8577, 8577, 8577, 8577, 8577,
  8971, 9072, 8964, 8965, 8965, 8966, 8967, 8967, 8967, 8968, 8968, 8968, 
    8968, 8968, 8968, 9066, 9002, 9002, 9002, 9002, 9002, 9002,
  8960, 9061, 8941, 8942, 8942, 8943, 8944, 8944, 8944, 8945, 8945, 8945, 
    8945, 8945, 8945, 9053, 8983, 8983, 8983, 8983, 8983, 8983,
  8922, 9019, 8763, 8760, 8758, 8756, 8756, 8755, 8754, 8750, 8750, 8750, 
    8750, 8750, 8750, 8886, 8653, 8653, 8653, 8653, 8653, 8653,
  8983, 9082, 8900, 8897, 8894, 8893, 8892, 8891, 8890, 8886, 8886, 8886, 
    8886, 8886, 8886, 8993, 8782, 8782, 8782, 8782, 8782, 8782,
  9009, 9109, 8771, 8765, 8760, 8756, 8754, 8752, 8749, 8742, 8742, 8742, 
    8742, 8742, 8742, 8913, 8505, 8505, 8505, 8505, 8505, 8505,
  8995, 9093, 8840, 8839, 8838, 8837, 8838, 8837, 8837, 8835, 8835, 8835, 
    8835, 8835, 8835, 8985, 8802, 8802, 8802, 8802, 8802, 8802,
  8921, 9020, 8794, 8791, 8790, 8788, 8788, 8787, 8787, 8784, 8784, 8784, 
    8784, 8784, 8784, 8919, 8710, 8710, 8710, 8710, 8710, 8710,
  9004, 9102, 8742, 8740, 8739, 8738, 8738, 8737, 8737, 8735, 8735, 8735, 
    8735, 8735, 8735, 8939, 8678, 8678, 8678, 8678, 8678, 8678,
  9092, 9187, 8738, 8737, 8736, 8735, 8735, 8735, 8734, 8732, 8732, 8732, 
    8732, 8732, 8732, 8973, 8689, 8689, 8689, 8689, 8689, 8689,
  9164, 9253, 8871, 8868, 8866, 8864, 8864, 8863, 8862, 8859, 8859, 8859, 
    8859, 8859, 8859, 9029, 8764, 8764, 8764, 8764, 8764, 8764,
  9105, 9195, 8891, 8887, 8885, 8884, 8883, 8882, 8881, 8877, 8877, 8877, 
    8877, 8877, 8877, 9015, 8772, 8772, 8772, 8772, 8772, 8772,
  9167, 9252, 8876, 8872, 8869, 8867, 8866, 8864, 8863, 8858, 8858, 8858, 
    8858, 8858, 8858, 9005, 8714, 8714, 8714, 8714, 8714, 8714,
  9265, 9347, 8912, 8908, 8906, 8905, 8904, 8903, 8902, 8898, 8898, 8898, 
    8898, 8898, 8898, 9069, 8788, 8788, 8788, 8788, 8788, 8788,
  9374, 9452, 9006, 9003, 9001, 8999, 8998, 8997, 8995, 8992, 8992, 8992, 
    8992, 8992, 8992, 9151, 8872, 8872, 8872, 8872, 8872, 8872,
  9314, 9395, 8972, 8969, 8966, 8964, 8963, 8962, 8960, 8956, 8956, 8956, 
    8956, 8956, 8956, 9112, 8827, 8827, 8827, 8827, 8827, 8827,
  9282, 9365, 8958, 8955, 8953, 8952, 8951, 8950, 8949, 8946, 8946, 8946, 
    8946, 8946, 8946, 9106, 8849, 8849, 8849, 8849, 8849, 8849,
  9173, 9262, 8936, 8933, 8932, 8930, 8930, 8929, 8928, 8925, 8925, 8925, 
    8925, 8925, 8925, 9069, 8843, 8843, 8843, 8843, 8843, 8843,
  8994, 9092, 8785, 8784, 8783, 8783, 8783, 8783, 8782, 8781, 8781, 8781, 
    8781, 8781, 8781, 8958, 8753, 8753, 8753, 8753, 8753, 8753,
  8774, 8883, 8636, 8637, 8637, 8637, 8638, 8638, 8639, 8639, 8639, 8639, 
    8639, 8639, 8639, 8839, 8666, 8666, 8666, 8666, 8666, 8666,
  8674, 8789, 8569, 8570, 8571, 8572, 8574, 8574, 8575, 8576, 8576, 8576, 
    8576, 8576, 8576, 8785, 8633, 8633, 8633, 8633, 8633, 8633,
  8172, 8317, 8130, 8135, 8139, 8142, 8147, 8149, 8151, 8157, 8157, 8157, 
    8157, 8157, 8157, 8493, 8384, 8384, 8384, 8384, 8384, 8384,
  8225, 8366, 8109, 8115, 8119, 8122, 8127, 8129, 8131, 8137, 8137, 8137, 
    8137, 8137, 8137, 8495, 8370, 8370, 8370, 8370, 8370, 8370,
  8160, 8303, 8267, 8273, 8277, 8280, 8285, 8287, 8289, 8296, 8296, 8296, 
    8296, 8296, 8296, 8554, 8540, 8540, 8540, 8540, 8540, 8540,
  8209, 8349, 8281, 8286, 8290, 8293, 8297, 8299, 8301, 8308, 8308, 8308, 
    8308, 8308, 8308, 8564, 8531, 8531, 8531, 8531, 8531, 8531,
  8207, 8348, 7962, 7969, 7973, 7977, 7981, 7983, 7986, 7993, 7993, 7993, 
    7993, 7993, 7993, 8420, 8243, 8243, 8243, 8243, 8243, 8243,
  8242, 8381, 8028, 8034, 8038, 8041, 8045, 8048, 8050, 8056, 8056, 8056, 
    8056, 8056, 8056, 8460, 8289, 8289, 8289, 8289, 8289, 8289,
  8293, 8426, 8154, 8158, 8160, 8162, 8166, 8167, 8168, 8173, 8173, 8173, 
    8173, 8173, 8173, 8496, 8334, 8334, 8334, 8334, 8334, 8334,
  8165, 8303, 8074, 8078, 8080, 8083, 8086, 8087, 8089, 8093, 8093, 8093, 
    8093, 8093, 8093, 8408, 8255, 8255, 8255, 8255, 8255, 8255,
  8018, 8154, 7861, 7864, 7867, 7869, 7872, 7874, 7875, 7879, 7879, 7879, 
    7879, 7879, 7879, 8214, 8032, 8032, 8032, 8032, 8032, 8032,
  7997, 8148, 8060, 8069, 8075, 8080, 8086, 8089, 8093, 8103, 8103, 8103, 
    8103, 8103, 8103, 8431, 8458, 8458, 8458, 8458, 8458, 8458,
  7991, 8142, 8081, 8089, 8096, 8100, 8106, 8109, 8112, 8121, 8121, 8121, 
    8121, 8121, 8121, 8431, 8456, 8456, 8456, 8456, 8456, 8456,
  8140, 8276, 8014, 8004, 7997, 7992, 7988, 7985, 7981, 7970, 7970, 7970, 
    7970, 7970, 7970, 8210, 7611, 7611, 7611, 7611, 7611, 7611,
  8126, 8268, 8206, 8212, 8217, 8220, 8225, 8227, 8229, 8236, 8236, 8236, 
    8236, 8236, 8236, 8501, 8488, 8488, 8488, 8488, 8488, 8488,
  8282, 8416, 8290, 8295, 8299, 8302, 8305, 8307, 8309, 8315, 8315, 8315, 
    8315, 8315, 8315, 8572, 8521, 8521, 8521, 8521, 8521, 8521,
  8241, 8377, 8304, 8309, 8313, 8316, 8320, 8322, 8324, 8330, 8330, 8330, 
    8330, 8330, 8330, 8569, 8547, 8547, 8547, 8547, 8547, 8547,
  8297, 8421, 8099, 8099, 8099, 8098, 8099, 8099, 8099, 8099, 8099, 8099, 
    8099, 8099, 8099, 8377, 8099, 8099, 8099, 8099, 8099, 8099,
  8277, 8407, 8029, 8030, 8031, 8031, 8033, 8033, 8034, 8035, 8035, 8035, 
    8035, 8035, 8035, 8382, 8088, 8088, 8088, 8088, 8088, 8088,
  8156, 8296, 8182, 8187, 8191, 8194, 8198, 8200, 8202, 8208, 8208, 8208, 
    8208, 8208, 8208, 8490, 8428, 8428, 8428, 8428, 8428, 8428,
  8230, 8382, 8147, 8155, 8161, 8165, 8170, 8173, 8176, 8185, 8185, 8185, 
    8185, 8185, 8185, 8595, 8499, 8499, 8499, 8499, 8499, 8499,
  8160, 8312, 7929, 7940, 7948, 7954, 7961, 7965, 7969, 7982, 7982, 7982, 
    7982, 7982, 7982, 8491, 8423, 8423, 8423, 8423, 8423, 8423,
  7895, 8059, 7693, 7707, 7717, 7724, 7732, 7737, 7742, 7757, 7757, 7757, 
    7757, 7757, 7757, 8307, 8280, 8280, 8280, 8280, 8280, 8280,
  7503, 7686, 7447, 7466, 7480, 7491, 7502, 7509, 7516, 7537, 7537, 7537, 
    7537, 7537, 7537, 8132, 8278, 8278, 8278, 8278, 8278, 8278,
  7295, 7489, 7270, 7290, 7304, 7314, 7326, 7333, 7340, 7362, 7362, 7362, 
    7362, 7362, 7362, 7990, 8117, 8117, 8117, 8117, 8117, 8117,
  6986, 7205, 6964, 6986, 7001, 7013, 7026, 7034, 7041, 7066, 7066, 7066, 
    7066, 7066, 7066, 7817, 7898, 7898, 7898, 7898, 7898, 7898,
  6553, 6797, 6524, 6552, 6571, 6586, 6602, 6612, 6621, 6652, 6652, 6652, 
    6652, 6652, 6652, 7552, 7699, 7699, 7698, 7698, 7698, 7698,
  6320, 6577, 6005, 6040, 6064, 6083, 6103, 6116, 6128, 6167, 6167, 6167, 
    6167, 6167, 6167, 7315, 7497, 7497, 7497, 7497, 7497, 7497,
  6038, 6256, 6078, 6106, 6127, 6142, 6157, 6167, 6178, 6211, 6211, 6211, 
    6211, 6211, 6211, 7318, 7469, 7607, 7607, 7607, 7607, 7607,
  6040, 6241, 5887, 5914, 5933, 5949, 5963, 5972, 5983, 6015, 6015, 6015, 
    6015, 6015, 6015, 7273, 7292, 7435, 7435, 7435, 7435, 7435,
  6108, 6293, 5904, 5929, 5948, 5962, 5975, 5984, 5995, 6025, 6025, 6025, 
    6025, 6025, 6025, 7266, 7259, 7400, 7400, 7400, 7400, 7400,
  6630, 6796, 6061, 6104, 6135, 6158, 6180, 6195, 6210, 6258, 6258, 6258, 
    6258, 6258, 6258, 7583, 7869, 7869, 7869, 7869, 7869, 7869,
  6638, 6769, 5943, 5988, 6020, 6043, 6067, 6082, 6098, 6147, 6147, 6147, 
    6147, 6147, 6147, 7476, 7814, 7814, 7814, 7814, 7813, 7814,
  6497, 6679, 6258, 6282, 6299, 6312, 6325, 6333, 6343, 6371, 6371, 6371, 
    6371, 6371, 6371, 7585, 7505, 7638, 7638, 7638, 7638, 7638,
  6639, 6849, 6668, 6693, 6711, 6725, 6738, 6746, 6756, 6785, 6785, 6785, 
    6785, 6785, 6785, 7783, 7859, 7980, 7980, 7980, 7980, 7980,
  6634, 6859, 6824, 6850, 6869, 6883, 6896, 6905, 6916, 6945, 6945, 6945, 
    6945, 6945, 6945, 7823, 8006, 8123, 8123, 8123, 8123, 8123,
  6540, 6785, 6849, 6877, 6897, 6912, 6927, 6936, 6948, 6980, 6980, 6980, 
    6980, 6980, 6980, 7817, 8079, 8197, 8197, 8197, 8197, 8197,
  6363, 6600, 6665, 6693, 6713, 6729, 6743, 6753, 6764, 6796, 6796, 6796, 
    6796, 6796, 6796, 7630, 7923, 8044, 8044, 8044, 8044, 8044,
  6150, 6396, 6398, 6428, 6449, 6465, 6481, 6491, 6503, 6537, 6537, 6537, 
    6537, 6537, 6537, 7498, 7761, 7890, 7890, 7890, 7890, 7890,
  5924, 6170, 6025, 6057, 6079, 6096, 6113, 6124, 6136, 6172, 6172, 6172, 
    6172, 6172, 6172, 7332, 7505, 7645, 7645, 7645, 7645, 7645,
  6004, 6217, 5712, 5764, 5801, 5828, 5855, 5872, 5891, 5948, 5948, 5948, 
    5948, 5948, 5948, 7254, 7870, 7870, 7870, 7870, 7870, 7870,
  5826, 6044, 5515, 5568, 5606, 5634, 5662, 5680, 5699, 5757, 5757, 5757, 
    5757, 5757, 5757, 7124, 7734, 7733, 7734, 7734, 7733, 7734,
  5391, 5624, 5306, 5339, 5362, 5381, 5398, 5409, 5422, 5461, 5461, 5461, 
    5461, 5461, 5461, 6853, 6967, 7127, 7127, 7127, 7127, 7127,
  5202, 5456, 5187, 5223, 5248, 5268, 5286, 5299, 5313, 5355, 5355, 5355, 
    5355, 5355, 5355, 6780, 6944, 7107, 7107, 7107, 7107, 7107,
  5031, 5306, 5136, 5174, 5201, 5222, 5242, 5255, 5270, 5314, 5314, 5314, 
    5314, 5314, 5314, 6709, 6961, 7127, 7127, 7127, 7127, 7127,
  4948, 5231, 5173, 5212, 5240, 5261, 5281, 5295, 5310, 5355, 5355, 5355, 
    5355, 5355, 5355, 6659, 7006, 7170, 7170, 7170, 7170, 7170,
  4928, 5211, 5166, 5205, 5232, 5254, 5274, 5288, 5303, 5348, 5348, 5348, 
    5348, 5348, 5348, 6642, 7002, 7166, 7166, 7166, 7166, 7166,
  5005, 5288, 5223, 5262, 5290, 5311, 5331, 5345, 5359, 5404, 5404, 5404, 
    5404, 5404, 5404, 6708, 7043, 7206, 7206, 7206, 7206, 7206,
  5302, 5577, 5535, 5572, 5598, 5618, 5637, 5650, 5664, 5706, 5706, 5706, 
    5706, 5706, 5706, 6920, 7240, 7395, 7395, 7395, 7395, 7395,
  5712, 5954, 6092, 6123, 6145, 6162, 6178, 6189, 6201, 6237, 6237, 6237, 
    6237, 6237, 6237, 7098, 7533, 7668, 7668, 7668, 7668, 7668,
  6341, 6588, 6903, 6931, 6952, 6967, 6982, 6991, 7002, 7034, 7034, 7034, 
    7034, 7034, 7034, 7617, 8110, 8224, 8224, 8224, 8224, 8224,
  6906, 7162, 7608, 7634, 7653, 7667, 7680, 7689, 7700, 7729, 7729, 7729, 
    7729, 7729, 7729, 8110, 8625, 8720, 8720, 8720, 8720, 8720,
  7360, 7691, 7896, 7907, 7915, 7921, 7927, 7930, 7934, 7946, 7946, 7946, 
    7946, 7946, 7946, 8406, 8357, 8357, 8357, 8357, 8357, 8357,
  7584, 7766, 7681, 7696, 7706, 7713, 7720, 7724, 7729, 7745, 7745, 7745, 
    7745, 7745, 7745, 8074, 8262, 8262, 8262, 8262, 8262, 8262,
  7946, 8093, 7791, 7800, 7807, 7812, 7819, 7822, 7825, 7836, 7836, 7836, 
    7836, 7836, 7836, 8260, 8210, 8210, 8210, 8210, 8210, 8210,
  7987, 8130, 8038, 8046, 8052, 8056, 8062, 8065, 8068, 8077, 8077, 8077, 
    8077, 8077, 8077, 8367, 8397, 8397, 8397, 8397, 8397, 8397,
  8042, 8189, 8427, 8431, 8434, 8437, 8440, 8441, 8443, 8448, 8448, 8448, 
    8448, 8448, 8448, 8564, 8618, 8618, 8618, 8618, 8618, 8618,
  7878, 8192, 8503, 8494, 8487, 8482, 8477, 8474, 8470, 8460, 8460, 8460, 
    8460, 8460, 8460, 8519, 8101, 8101, 8101, 8101, 8101, 8101,
  7756, 7901, 8288, 8300, 8309, 8316, 8322, 8326, 8331, 8345, 8345, 8345, 
    8345, 8345, 8345, 8363, 8799, 8869, 8869, 8869, 8869, 8869,
  7298, 7641, 8057, 8054, 8052, 8050, 8048, 8047, 8045, 8042, 8042, 8042, 
    8042, 8042, 8042, 8144, 7915, 7915, 7915, 7915, 7915, 7915,
  6948, 7220, 7571, 7569, 7568, 7567, 7566, 7565, 7564, 7562, 7562, 7562, 
    7562, 7562, 7562, 7519, 7489, 7489, 7489, 7489, 7489, 7490,
  6567, 6916, 7470, 7467, 7465, 7463, 7462, 7460, 7459, 7455, 7455, 7455, 
    7455, 7455, 7455, 7416, 7333, 7333, 7333, 7333, 7333, 7333,
  6326, 6785, 7580, 7576, 7573, 7570, 7567, 7565, 7563, 7558, 7558, 7558, 
    7558, 7558, 7558, 7589, 7373, 7373, 7372, 7372, 7373, 7373,
  8680, 8790, 8905, 8909, 8912, 8914, 8917, 8918, 8919, 8923, 8923, 8923, 
    8923, 8923, 8923, 8955, 9074, 9074, 9074, 9074, 9074, 9074,
  8745, 8853, 8931, 8932, 8933, 8934, 8936, 8936, 8937, 8939, 8939, 8939, 
    8939, 8939, 8939, 8974, 9008, 9008, 9008, 9008, 9008, 9008,
  8817, 8924, 8961, 8961, 8962, 8962, 8963, 8963, 8964, 8964, 8964, 8964, 
    8964, 8964, 8964, 9012, 8995, 8995, 8995, 8995, 8995, 8995,
  8911, 9016, 9054, 9056, 9058, 9059, 9061, 9062, 9063, 9066, 9066, 9066, 
    9066, 9066, 9066, 9118, 9170, 9170, 9170, 9170, 9170, 9170,
  8963, 9063, 9083, 9084, 9086, 9086, 9088, 9089, 9089, 9091, 9091, 9091, 
    9091, 9091, 9091, 9127, 9164, 9164, 9164, 9164, 9164, 9164,
  9041, 9133, 9131, 9137, 9141, 9144, 9148, 9150, 9152, 9158, 9158, 9158, 
    9158, 9158, 9158, 9195, 9384, 9384, 9384, 9384, 9384, 9384,
  8965, 9064, 9026, 9029, 9031, 9033, 9035, 9036, 9037, 9041, 9041, 9041, 
    9041, 9041, 9041, 9110, 9159, 9159, 9159, 9159, 9159, 9159,
  8898, 9005, 8950, 8952, 8954, 8955, 8957, 8958, 8958, 8961, 8961, 8961, 
    8961, 8961, 8961, 9065, 9049, 9049, 9049, 9049, 9049, 9049,
  8858, 8965, 8910, 8914, 8918, 8920, 8924, 8925, 8927, 8932, 8932, 8932, 
    8932, 8932, 8932, 9049, 9120, 9120, 9120, 9120, 9120, 9120,
  8841, 8951, 8902, 8903, 8903, 8903, 8905, 8905, 8905, 8906, 8906, 8906, 
    8906, 8906, 8906, 9007, 8935, 8935, 8935, 8935, 8935, 8935,
  8959, 9061, 8965, 8964, 8964, 8963, 8964, 8963, 8963, 8962, 8962, 8962, 
    8962, 8962, 8962, 9047, 8934, 8934, 8934, 8934, 8934, 8934,
  9034, 9127, 8994, 8990, 8988, 8986, 8985, 8984, 8982, 8979, 8979, 8979, 
    8979, 8979, 8979, 9033, 8858, 8858, 8858, 8858, 8858, 8858,
  8867, 8961, 8753, 8748, 8744, 8741, 8740, 8738, 8736, 8730, 8730, 8730, 
    8730, 8730, 8730, 8808, 8547, 8547, 8547, 8547, 8547, 8547,
  9133, 9201, 8993, 8980, 8970, 8963, 8957, 8953, 8948, 8933, 8933, 8933, 
    8933, 8933, 8933, 8858, 8448, 8448, 8448, 8448, 8448, 8448,
  8963, 9046, 8753, 8743, 8737, 8731, 8727, 8724, 8720, 8709, 8709, 8709, 
    8709, 8709, 8709, 8760, 8354, 8354, 8354, 8354, 8354, 8354,
  9076, 9167, 8964, 8963, 8963, 8962, 8963, 8962, 8962, 8961, 8961, 8961, 
    8961, 8961, 8961, 9063, 8942, 8942, 8942, 8942, 8942, 8942,
  8891, 8996, 8879, 8881, 8882, 8882, 8884, 8884, 8885, 8886, 8886, 8886, 
    8886, 8886, 8886, 9007, 8941, 8941, 8941, 8941, 8941, 8941,
  8833, 8938, 8609, 8609, 8608, 8608, 8609, 8609, 8609, 8608, 8608, 8608, 
    8608, 8608, 8608, 8827, 8602, 8602, 8602, 8602, 8602, 8602,
  8970, 9070, 8832, 8831, 8831, 8831, 8832, 8832, 8832, 8831, 8831, 8831, 
    8831, 8831, 8831, 8991, 8831, 8831, 8831, 8831, 8831, 8831,
  8953, 9054, 8801, 8802, 8802, 8802, 8803, 8804, 8804, 8804, 8804, 8804, 
    8804, 8804, 8804, 8978, 8828, 8828, 8828, 8828, 8828, 8828,
  8967, 9067, 8808, 8808, 8808, 8807, 8808, 8808, 8808, 8808, 8808, 8808, 
    8808, 8808, 8808, 8974, 8811, 8811, 8811, 8811, 8811, 8811,
  8932, 9033, 8758, 8757, 8755, 8754, 8754, 8754, 8753, 8751, 8751, 8751, 
    8751, 8751, 8751, 8920, 8694, 8694, 8694, 8694, 8694, 8694,
  8895, 9002, 8578, 8580, 8581, 8581, 8583, 8584, 8584, 8586, 8586, 8586, 
    8586, 8586, 8586, 8878, 8648, 8648, 8648, 8648, 8648, 8648,
  9045, 9144, 8713, 8714, 8714, 8714, 8715, 8716, 8716, 8716, 8716, 8716, 
    8716, 8716, 8716, 8973, 8741, 8741, 8741, 8741, 8741, 8741,
  9029, 9127, 8712, 8712, 8712, 8713, 8714, 8714, 8714, 8714, 8714, 8714, 
    8714, 8714, 8714, 8956, 8734, 8734, 8734, 8734, 8734, 8734,
  9093, 9184, 8817, 8815, 8814, 8813, 8813, 8812, 8812, 8810, 8810, 8810, 
    8810, 8810, 8810, 8987, 8749, 8749, 8749, 8749, 8749, 8749,
  9256, 9339, 8986, 8982, 8979, 8977, 8975, 8974, 8973, 8968, 8968, 8968, 
    8968, 8968, 8968, 9093, 8823, 8823, 8823, 8823, 8823, 8823,
  9351, 9427, 9013, 9010, 9008, 9006, 9005, 9004, 9003, 8999, 8999, 8999, 
    8999, 8999, 8999, 9137, 8889, 8889, 8889, 8889, 8889, 8889,
  9331, 9412, 8976, 8973, 8971, 8970, 8969, 8968, 8967, 8964, 8964, 8964, 
    8964, 8964, 8964, 9134, 8866, 8866, 8866, 8866, 8866, 8866,
  9504, 9582, 9274, 9264, 9257, 9252, 9248, 9245, 9241, 9230, 9230, 9230, 
    9230, 9230, 9230, 9286, 8875, 8875, 8875, 8875, 8875, 8875,
  9270, 9352, 8989, 8986, 8984, 8982, 8981, 8980, 8979, 8975, 8975, 8975, 
    8975, 8975, 8975, 9108, 8865, 8865, 8866, 8866, 8865, 8865,
  9125, 9214, 8909, 8907, 8905, 8904, 8904, 8903, 8902, 8900, 8900, 8900, 
    8900, 8900, 8900, 9038, 8826, 8826, 8826, 8826, 8826, 8826,
  8900, 9001, 8739, 8738, 8737, 8737, 8737, 8737, 8737, 8736, 8736, 8736, 
    8736, 8736, 8736, 8901, 8717, 8717, 8717, 8717, 8717, 8717,
  8982, 9079, 8770, 8770, 8769, 8769, 8770, 8770, 8769, 8769, 8769, 8769, 
    8769, 8769, 8769, 8944, 8759, 8759, 8759, 8759, 8759, 8759,
  8551, 8673, 8447, 8449, 8450, 8452, 8454, 8455, 8455, 8458, 8458, 8458, 
    8458, 8458, 8458, 8707, 8549, 8549, 8549, 8549, 8549, 8549,
  8208, 8348, 8141, 8146, 8149, 8152, 8156, 8158, 8159, 8165, 8165, 8165, 
    8165, 8165, 8165, 8485, 8366, 8366, 8366, 8366, 8366, 8366,
  8008, 8162, 8194, 8201, 8206, 8209, 8214, 8216, 8219, 8226, 8226, 8226, 
    8226, 8226, 8226, 8490, 8496, 8496, 8496, 8496, 8496, 8496,
  7887, 8046, 7772, 7781, 7788, 7793, 7799, 7802, 7805, 7815, 7815, 7815, 
    7815, 7815, 7815, 8274, 8167, 8167, 8167, 8167, 8167, 8167,
  7952, 8105, 7801, 7809, 7814, 7818, 7823, 7826, 7828, 7837, 7837, 7837, 
    7837, 7837, 7837, 8272, 8129, 8129, 8129, 8129, 8129, 8129,
  8138, 8277, 7928, 7934, 7939, 7942, 7946, 7948, 7950, 7957, 7957, 7957, 
    7957, 7957, 7957, 8353, 8193, 8193, 8193, 8193, 8193, 8193,
  8316, 8445, 8138, 8141, 8144, 8146, 8149, 8151, 8152, 8156, 8156, 8156, 
    8156, 8156, 8156, 8478, 8308, 8308, 8308, 8308, 8308, 8308,
  8359, 8490, 8123, 8127, 8130, 8132, 8136, 8137, 8139, 8143, 8143, 8143, 
    8143, 8143, 8143, 8509, 8310, 8310, 8310, 8310, 8310, 8310,
  8218, 8358, 7963, 7966, 7967, 7968, 7971, 7972, 7972, 7975, 7975, 7975, 
    7975, 7975, 7975, 8382, 8073, 8073, 8073, 8073, 8073, 8073,
  8080, 8223, 7899, 7904, 7908, 7911, 7915, 7917, 7918, 7924, 7924, 7924, 
    7924, 7924, 7924, 8319, 8133, 8133, 8133, 8133, 8133, 8133,
  8172, 8317, 7982, 7982, 7982, 7981, 7982, 7982, 7982, 7981, 7981, 7981, 
    7981, 7981, 7981, 8358, 7977, 7977, 7977, 7977, 7977, 7977,
  8148, 8289, 8155, 8161, 8165, 8169, 8173, 8175, 8177, 8184, 8184, 8184, 
    8184, 8184, 8184, 8478, 8420, 8420, 8420, 8420, 8420, 8420,
  8138, 8280, 8167, 8173, 8177, 8180, 8185, 8187, 8189, 8196, 8196, 8196, 
    8196, 8196, 8196, 8483, 8436, 8436, 8436, 8436, 8436, 8436,
  8167, 8308, 8205, 8211, 8216, 8219, 8223, 8225, 8227, 8234, 8234, 8234, 
    8234, 8234, 8234, 8509, 8471, 8471, 8471, 8471, 8471, 8471,
  8188, 8327, 8239, 8245, 8248, 8251, 8255, 8257, 8259, 8266, 8266, 8266, 
    8266, 8266, 8266, 8526, 8485, 8485, 8485, 8485, 8485, 8485,
  8265, 8396, 8103, 8104, 8104, 8104, 8106, 8106, 8106, 8106, 8106, 8106, 
    8106, 8106, 8106, 8410, 8135, 8135, 8135, 8135, 8135, 8135,
  8262, 8393, 8126, 8127, 8128, 8129, 8131, 8131, 8132, 8133, 8133, 8133, 
    8133, 8133, 8133, 8429, 8192, 8192, 8192, 8192, 8192, 8192,
  8248, 8384, 8272, 8277, 8281, 8284, 8287, 8289, 8291, 8296, 8296, 8296, 
    8296, 8296, 8296, 8555, 8495, 8495, 8495, 8495, 8495, 8495,
  8228, 8365, 8255, 8260, 8263, 8266, 8269, 8271, 8273, 8278, 8278, 8278, 
    8278, 8278, 8278, 8540, 8474, 8474, 8474, 8474, 8474, 8474,
  8378, 8526, 8369, 8370, 8370, 8371, 8372, 8373, 8373, 8374, 8374, 8374, 
    8374, 8374, 8374, 8686, 8421, 8421, 8421, 8421, 8421, 8421,
  8136, 8281, 8242, 8246, 8249, 8251, 8255, 8256, 8258, 8263, 8263, 8263, 
    8263, 8263, 8263, 8518, 8436, 8436, 8436, 8436, 8436, 8436,
  7936, 8095, 7991, 7997, 8001, 8005, 8009, 8011, 8013, 8020, 8020, 8020, 
    8020, 8020, 8020, 8370, 8259, 8259, 8259, 8259, 8259, 8259,
  7643, 7821, 7614, 7630, 7641, 7650, 7659, 7665, 7670, 7688, 7688, 7688, 
    7688, 7688, 7688, 8227, 8292, 8292, 8292, 8292, 8292, 8292,
  7313, 7508, 7283, 7302, 7315, 7325, 7336, 7343, 7349, 7370, 7370, 7370, 
    7370, 7370, 7370, 8001, 8090, 8090, 8090, 8090, 8090, 8090,
  6819, 7043, 6566, 6596, 6617, 6633, 6649, 6660, 6670, 6704, 6704, 6704, 
    6704, 6704, 6704, 7641, 7826, 7826, 7826, 7826, 7826, 7826,
  6506, 6757, 6065, 6099, 6122, 6141, 6160, 6172, 6183, 6221, 6221, 6221, 
    6221, 6221, 6221, 7400, 7497, 7497, 7497, 7497, 7497, 7497,
  5801, 6028, 5811, 5841, 5863, 5880, 5896, 5906, 5918, 5954, 5954, 5954, 
    5954, 5954, 5954, 7160, 7306, 7452, 7452, 7452, 7452, 7452,
  5466, 5714, 5555, 5588, 5612, 5631, 5648, 5660, 5673, 5713, 5713, 5713, 
    5713, 5713, 5713, 6963, 7186, 7339, 7339, 7339, 7339, 7339,
  5382, 5646, 5604, 5639, 5664, 5684, 5702, 5714, 5728, 5769, 5769, 5769, 
    5769, 5769, 5769, 6940, 7257, 7409, 7409, 7409, 7409, 7409,
  5425, 5681, 5685, 5719, 5744, 5762, 5780, 5792, 5805, 5845, 5845, 5845, 
    5845, 5845, 5845, 6937, 7292, 7441, 7441, 7441, 7441, 7441,
  5611, 5854, 5730, 5762, 5786, 5803, 5820, 5832, 5844, 5882, 5882, 5882, 
    5882, 5882, 5882, 7056, 7290, 7438, 7438, 7438, 7438, 7438,
  5835, 6051, 5827, 5856, 5877, 5893, 5908, 5918, 5930, 5964, 5964, 5964, 
    5964, 5964, 5964, 7142, 7287, 7431, 7431, 7431, 7431, 7431,
  6140, 6353, 6210, 6237, 6257, 6272, 6286, 6296, 6307, 6338, 6338, 6338, 
    6338, 6338, 6338, 7378, 7551, 7685, 7685, 7685, 7685, 7685,
  6381, 6616, 6626, 6654, 6674, 6689, 6704, 6713, 6724, 6756, 6756, 6756, 
    6756, 6756, 6756, 7648, 7896, 8019, 8019, 8019, 8019, 8019,
  6538, 6760, 6823, 6849, 6868, 6882, 6895, 6904, 6914, 6944, 6944, 6944, 
    6944, 6944, 6944, 7713, 7990, 8107, 8107, 8107, 8107, 8107,
  6602, 6844, 6930, 6957, 6977, 6992, 7006, 7015, 7026, 7057, 7057, 7057, 
    7057, 7057, 7057, 7848, 8123, 8237, 8237, 8237, 8237, 8237,
  6563, 6809, 6850, 6878, 6898, 6913, 6928, 6937, 6949, 6980, 6980, 6980, 
    6980, 6980, 6980, 7839, 8080, 8197, 8197, 8197, 8197, 8197,
  6424, 6664, 6595, 6624, 6644, 6660, 6674, 6684, 6695, 6728, 6728, 6728, 
    6728, 6728, 6728, 7711, 7883, 8007, 8007, 8007, 8007, 8007,
  6227, 6474, 6363, 6393, 6415, 6431, 6447, 6457, 6469, 6504, 6504, 6504, 
    6504, 6504, 6504, 7587, 7747, 7879, 7879, 7879, 7879, 7879,
  5975, 6195, 5978, 6007, 6028, 6044, 6059, 6069, 6080, 6114, 6114, 6114, 
    6114, 6114, 6114, 7276, 7404, 7544, 7544, 7544, 7544, 7544,
  5774, 6016, 5821, 5853, 5876, 5893, 5910, 5921, 5933, 5970, 5970, 5970, 
    5970, 5970, 5970, 7196, 7350, 7496, 7496, 7496, 7496, 7496,
  5556, 5806, 5583, 5617, 5641, 5659, 5677, 5688, 5701, 5741, 5741, 5741, 
    5741, 5741, 5741, 7054, 7209, 7362, 7362, 7362, 7362, 7362,
  5284, 5537, 5313, 5348, 5373, 5393, 5411, 5423, 5437, 5478, 5478, 5478, 
    5478, 5478, 5478, 6841, 7030, 7190, 7190, 7190, 7190, 7190,
  5066, 5341, 5188, 5226, 5252, 5273, 5293, 5306, 5321, 5365, 5365, 5365, 
    5365, 5365, 5365, 6736, 6997, 7162, 7162, 7162, 7162, 7162,
  4895, 5176, 5129, 5168, 5196, 5217, 5237, 5251, 5266, 5311, 5311, 5311, 
    5311, 5311, 5311, 6601, 6966, 7131, 7131, 7131, 7131, 7131,
  4845, 5126, 5058, 5097, 5125, 5146, 5167, 5181, 5195, 5241, 5241, 5241, 
    5241, 5241, 5241, 6563, 6917, 7083, 7083, 7083, 7083, 7083,
  4987, 5266, 5207, 5246, 5273, 5294, 5314, 5327, 5342, 5386, 5386, 5386, 
    5386, 5386, 5386, 6673, 7018, 7181, 7181, 7181, 7181, 7181,
  5328, 5603, 5555, 5591, 5617, 5637, 5656, 5669, 5683, 5725, 5725, 5725, 
    5725, 5725, 5725, 6941, 7254, 7408, 7408, 7408, 7408, 7408,
  5848, 6093, 6120, 6152, 6174, 6191, 6207, 6218, 6230, 6266, 6266, 6266, 
    6266, 6266, 6266, 7239, 7563, 7699, 7699, 7699, 7699, 7699,
  6439, 6656, 6881, 6907, 6925, 6938, 6952, 6960, 6970, 6999, 6999, 6999, 
    6999, 6999, 6999, 7586, 8016, 8129, 8129, 8129, 8129, 8129,
  7117, 7455, 7704, 7723, 7736, 7745, 7754, 7760, 7766, 7787, 7787, 7787, 
    7787, 7787, 7787, 8292, 8455, 8455, 8455, 8455, 8455, 8455,
  7578, 7866, 7984, 7993, 7999, 8004, 8009, 8011, 8014, 8024, 8024, 8024, 
    8024, 8024, 8024, 8418, 8354, 8354, 8354, 8354, 8355, 8354,
  7834, 8046, 7996, 8004, 8010, 8014, 8018, 8020, 8023, 8032, 8032, 8032, 
    8032, 8032, 8032, 8353, 8325, 8325, 8325, 8325, 8325, 8325,
  8018, 8178, 8055, 8061, 8065, 8068, 8071, 8073, 8075, 8081, 8081, 8081, 
    8081, 8081, 8081, 8299, 8298, 8298, 8298, 8298, 8298, 8298,
  7997, 8144, 8195, 8206, 8213, 8219, 8225, 8229, 8232, 8244, 8244, 8244, 
    8244, 8244, 8244, 8491, 8644, 8644, 8644, 8644, 8644, 8644,
  7787, 7950, 8258, 8268, 8275, 8280, 8286, 8290, 8293, 8305, 8305, 8305, 
    8305, 8305, 8305, 8484, 8686, 8686, 8686, 8686, 8686, 8686,
  7835, 7998, 8391, 8397, 8401, 8404, 8408, 8410, 8412, 8419, 8419, 8419, 
    8419, 8419, 8419, 8529, 8650, 8650, 8650, 8650, 8650, 8650,
  7744, 7902, 8254, 8268, 8278, 8285, 8292, 8296, 8303, 8318, 8318, 8318, 
    8318, 8318, 8318, 8416, 8817, 8889, 8889, 8889, 8889, 8889,
  7612, 7773, 8092, 8106, 8117, 8125, 8132, 8137, 8143, 8159, 8159, 8159, 
    8159, 8159, 8159, 8317, 8707, 8784, 8784, 8784, 8784, 8784,
  7179, 7449, 7790, 7785, 7781, 7778, 7776, 7773, 7771, 7765, 7765, 7765, 
    7765, 7765, 7765, 7691, 7565, 7565, 7565, 7565, 7565, 7565,
  6720, 7050, 7576, 7570, 7566, 7562, 7559, 7556, 7554, 7546, 7546, 7546, 
    7546, 7546, 7546, 7443, 7300, 7300, 7300, 7300, 7300, 7300,
  6560, 7018, 7809, 7799, 7792, 7786, 7780, 7776, 7772, 7760, 7760, 7760, 
    7760, 7760, 7760, 7730, 7355, 7355, 7355, 7355, 7355, 7355,
  8730, 8838, 8990, 8992, 8994, 8995, 8997, 8997, 8998, 9001, 9001, 9001, 
    9001, 9001, 9001, 8999, 9094, 9094, 9094, 9094, 9094, 9094,
  8774, 8882, 9030, 9029, 9028, 9027, 9027, 9027, 9026, 9025, 9025, 9025, 
    9025, 9025, 9025, 9006, 8989, 8989, 8989, 8989, 8989, 8989,
  8874, 8978, 9050, 9049, 9048, 9047, 9048, 9047, 9047, 9045, 9045, 9045, 
    9045, 9045, 9045, 9052, 9010, 9010, 9010, 9010, 9010, 9010,
  8875, 8980, 9001, 9002, 9002, 9003, 9004, 9004, 9005, 9006, 9006, 9006, 
    9006, 9006, 9006, 9057, 9047, 9047, 9047, 9047, 9047, 9047,
  8945, 9046, 9121, 9122, 9122, 9123, 9124, 9125, 9125, 9126, 9126, 9126, 
    9126, 9126, 9126, 9130, 9175, 9175, 9175, 9175, 9175, 9175,
  8894, 8999, 8981, 8980, 8980, 8980, 8980, 8980, 8980, 8980, 8980, 8980, 
    8980, 8980, 8980, 9042, 8975, 8975, 8975, 8975, 8975, 8975,
  8945, 9044, 9062, 9067, 9070, 9072, 9076, 9077, 9079, 9085, 9085, 9085, 
    9085, 9085, 9085, 9133, 9272, 9272, 9272, 9272, 9272, 9272,
  8916, 9019, 9050, 9051, 9051, 9052, 9053, 9053, 9054, 9055, 9055, 9055, 
    9055, 9055, 9055, 9091, 9098, 9098, 9098, 9098, 9098, 9098,
  8986, 9089, 9031, 9030, 9030, 9029, 9030, 9029, 9029, 9028, 9028, 9028, 
    9028, 9028, 9028, 9103, 9004, 9004, 9004, 9004, 9004, 9004,
  8934, 9036, 8952, 8952, 8951, 8951, 8951, 8951, 8951, 8950, 8950, 8950, 
    8950, 8950, 8950, 9032, 8932, 8932, 8932, 8932, 8932, 8932,
  9040, 9121, 8972, 8958, 8948, 8941, 8935, 8930, 8925, 8910, 8910, 8910, 
    8910, 8910, 8910, 8855, 8405, 8405, 8405, 8405, 8405, 8405,
  9006, 9106, 9008, 9008, 9007, 9007, 9008, 9008, 9008, 9008, 9008, 9008, 
    9008, 9008, 9008, 9091, 9012, 9012, 9012, 9012, 9012, 9012,
  8990, 9090, 9022, 9023, 9024, 9025, 9026, 9027, 9027, 9028, 9028, 9028, 
    9028, 9028, 9028, 9108, 9080, 9080, 9080, 9080, 9080, 9080,
  9000, 9100, 9059, 9059, 9060, 9060, 9062, 9062, 9062, 9063, 9063, 9063, 
    9063, 9063, 9063, 9124, 9104, 9104, 9104, 9104, 9104, 9104,
  9009, 9106, 9040, 9039, 9038, 9038, 9039, 9038, 9038, 9037, 9037, 9037, 
    9037, 9037, 9037, 9090, 9019, 9019, 9019, 9019, 9019, 9019,
  8731, 8844, 8566, 8565, 8564, 8564, 8564, 8564, 8563, 8562, 8562, 8562, 
    8562, 8562, 8562, 8783, 8530, 8530, 8530, 8530, 8530, 8530,
  8879, 8984, 8892, 8893, 8894, 8894, 8896, 8896, 8896, 8897, 8897, 8897, 
    8897, 8897, 8897, 9006, 8939, 8939, 8939, 8939, 8939, 8939,
  8906, 9003, 8670, 8668, 8667, 8666, 8666, 8665, 8664, 8662, 8662, 8662, 
    8662, 8662, 8662, 8840, 8596, 8596, 8596, 8596, 8596, 8596,
  9050, 9143, 8856, 8846, 8840, 8834, 8830, 8827, 8823, 8812, 8812, 8812, 
    8812, 8812, 8812, 8910, 8459, 8459, 8459, 8459, 8459, 8459,
  9012, 9111, 8869, 8869, 8870, 8870, 8871, 8871, 8871, 8872, 8872, 8872, 
    8872, 8872, 8872, 9036, 8902, 8902, 8902, 8902, 8902, 8902,
  8990, 9086, 8730, 8729, 8728, 8727, 8727, 8726, 8726, 8724, 8724, 8724, 
    8724, 8724, 8724, 8916, 8674, 8674, 8674, 8674, 8674, 8674,
  8959, 9059, 8792, 8791, 8790, 8790, 8790, 8790, 8789, 8788, 8788, 8788, 
    8788, 8788, 8788, 8956, 8765, 8765, 8765, 8765, 8765, 8765,
  9029, 9126, 8776, 8776, 8776, 8775, 8776, 8776, 8776, 8775, 8775, 8775, 
    8775, 8775, 8775, 8977, 8766, 8766, 8766, 8766, 8766, 8766,
  9095, 9190, 8792, 8792, 8791, 8791, 8792, 8792, 8792, 8791, 8791, 8791, 
    8791, 8791, 8791, 9010, 8781, 8781, 8781, 8781, 8781, 8781,
  9019, 9119, 8730, 8730, 8731, 8731, 8732, 8732, 8732, 8732, 8732, 8732, 
    8732, 8732, 8732, 8970, 8751, 8751, 8751, 8751, 8751, 8751,
  9134, 9222, 8964, 8960, 8957, 8955, 8954, 8953, 8951, 8947, 8947, 8947, 
    8947, 8947, 8947, 9045, 8806, 8806, 8806, 8806, 8806, 8806,
  9195, 9282, 9024, 9020, 9017, 9015, 9014, 9013, 9012, 9008, 9008, 9008, 
    9008, 9008, 9008, 9103, 8880, 8880, 8880, 8880, 8880, 8880,
  9261, 9342, 8962, 8959, 8956, 8954, 8953, 8952, 8951, 8947, 8947, 8947, 
    8947, 8947, 8947, 9083, 8824, 8824, 8824, 8824, 8824, 8824,
  9327, 9407, 8976, 8973, 8971, 8969, 8968, 8967, 8966, 8962, 8962, 8962, 
    8962, 8962, 8962, 9126, 8854, 8854, 8854, 8854, 8854, 8854,
  9321, 9402, 8987, 8984, 8982, 8981, 8980, 8979, 8978, 8974, 8974, 8974, 
    8974, 8974, 8974, 9132, 8869, 8869, 8869, 8869, 8869, 8869,
  9277, 9358, 8948, 8946, 8944, 8943, 8943, 8942, 8942, 8939, 8939, 8939, 
    8939, 8939, 8939, 9099, 8868, 8868, 8868, 8868, 8868, 8868,
  9051, 9146, 8822, 8820, 8819, 8818, 8818, 8818, 8817, 8816, 8816, 8816, 
    8816, 8816, 8816, 8989, 8769, 8769, 8769, 8769, 8769, 8769,
  8841, 8949, 8646, 8647, 8648, 8648, 8649, 8650, 8650, 8651, 8651, 8651, 
    8651, 8651, 8651, 8878, 8688, 8688, 8688, 8688, 8688, 8688,
  8491, 8615, 8266, 8269, 8272, 8274, 8276, 8278, 8279, 8283, 8283, 8283, 
    8283, 8283, 8283, 8609, 8426, 8426, 8426, 8426, 8426, 8426,
  8267, 8405, 8168, 8174, 8177, 8180, 8184, 8186, 8188, 8194, 8194, 8194, 
    8194, 8194, 8194, 8527, 8406, 8406, 8406, 8406, 8406, 8406,
  8157, 8298, 8086, 8092, 8096, 8098, 8102, 8104, 8106, 8112, 8112, 8112, 
    8112, 8112, 8112, 8445, 8330, 8330, 8330, 8330, 8330, 8330,
  8022, 8174, 8165, 8172, 8177, 8180, 8185, 8188, 8190, 8198, 8198, 8198, 
    8198, 8198, 8198, 8478, 8470, 8470, 8470, 8470, 8470, 8470,
  8153, 8299, 7960, 7967, 7972, 7976, 7981, 7984, 7986, 7995, 7995, 7995, 
    7995, 7995, 7995, 8429, 8283, 8283, 8283, 8283, 8283, 8283,
  8330, 8459, 8246, 8249, 8251, 8253, 8255, 8256, 8257, 8261, 8261, 8261, 
    8261, 8261, 8261, 8530, 8380, 8380, 8380, 8380, 8380, 8380,
  8282, 8411, 8192, 8195, 8196, 8198, 8200, 8201, 8202, 8205, 8205, 8205, 
    8205, 8205, 8205, 8473, 8313, 8313, 8313, 8313, 8313, 8313,
  8322, 8449, 8157, 8159, 8161, 8162, 8165, 8166, 8166, 8169, 8169, 8169, 
    8169, 8169, 8169, 8467, 8275, 8275, 8275, 8275, 8275, 8275,
  8396, 8530, 8180, 8183, 8185, 8187, 8190, 8191, 8193, 8196, 8196, 8196, 
    8196, 8196, 8196, 8561, 8335, 8335, 8335, 8335, 8335, 8335,
  8313, 8451, 8064, 8070, 8074, 8077, 8081, 8083, 8085, 8091, 8091, 8091, 
    8091, 8091, 8091, 8506, 8313, 8313, 8313, 8313, 8313, 8313,
  8250, 8392, 8106, 8112, 8115, 8118, 8122, 8124, 8126, 8131, 8131, 8131, 
    8131, 8131, 8131, 8508, 8339, 8339, 8339, 8339, 8339, 8339,
  8185, 8329, 8062, 8066, 8069, 8071, 8074, 8076, 8077, 8081, 8081, 8081, 
    8081, 8081, 8081, 8446, 8245, 8245, 8245, 8245, 8245, 8245,
  8347, 8493, 8237, 8240, 8242, 8244, 8246, 8247, 8248, 8251, 8251, 8251, 
    8251, 8251, 8251, 8618, 8371, 8371, 8371, 8371, 8371, 8371,
  8455, 8600, 8305, 8307, 8309, 8310, 8312, 8313, 8314, 8317, 8317, 8317, 
    8317, 8317, 8317, 8698, 8418, 8418, 8418, 8418, 8418, 8418,
  8233, 8369, 8264, 8269, 8273, 8275, 8279, 8281, 8283, 8288, 8288, 8288, 
    8288, 8288, 8288, 8542, 8489, 8489, 8489, 8489, 8489, 8489,
  8219, 8356, 8268, 8273, 8277, 8280, 8284, 8285, 8287, 8293, 8293, 8293, 
    8293, 8293, 8293, 8546, 8506, 8506, 8506, 8506, 8506, 8506,
  8147, 8289, 8243, 8248, 8252, 8255, 8259, 8261, 8263, 8270, 8270, 8270, 
    8270, 8270, 8270, 8522, 8495, 8495, 8495, 8495, 8495, 8495,
  8313, 8445, 8190, 8188, 8186, 8185, 8185, 8184, 8183, 8180, 8180, 8180, 
    8180, 8180, 8180, 8449, 8101, 8101, 8101, 8101, 8101, 8101,
  8264, 8398, 8172, 8175, 8176, 8178, 8180, 8181, 8181, 8184, 8184, 8184, 
    8184, 8184, 8184, 8478, 8283, 8283, 8283, 8283, 8283, 8283,
  8515, 8657, 8509, 8510, 8510, 8511, 8512, 8512, 8512, 8513, 8513, 8513, 
    8513, 8513, 8513, 8802, 8551, 8551, 8551, 8551, 8551, 8551,
  8361, 8500, 8289, 8291, 8293, 8294, 8296, 8297, 8298, 8301, 8301, 8301, 
    8301, 8301, 8301, 8608, 8401, 8401, 8401, 8401, 8401, 8401,
  8203, 8352, 8157, 8164, 8170, 8174, 8179, 8182, 8184, 8193, 8193, 8193, 
    8193, 8193, 8193, 8569, 8491, 8491, 8491, 8491, 8491, 8491,
  8050, 8203, 8050, 8057, 8063, 8067, 8072, 8074, 8077, 8085, 8085, 8085, 
    8085, 8085, 8085, 8449, 8381, 8381, 8381, 8381, 8381, 8381,
  7783, 7951, 7826, 7841, 7851, 7859, 7868, 7873, 7878, 7894, 7894, 7894, 
    7894, 7894, 7894, 8343, 8453, 8453, 8453, 8453, 8453, 8453,
  7405, 7596, 7426, 7445, 7458, 7467, 7478, 7485, 7491, 7512, 7512, 7512, 
    7512, 7512, 7512, 8095, 8214, 8214, 8214, 8214, 8214, 8214,
  7076, 7293, 6770, 6797, 6816, 6830, 6845, 6854, 6863, 6893, 6893, 6893, 
    6893, 6893, 6893, 7810, 7894, 7894, 7894, 7894, 7894, 7894,
  6424, 6534, 5817, 5864, 5897, 5921, 5946, 5961, 5978, 6030, 6030, 6030, 
    6030, 6030, 6030, 7188, 7765, 7764, 7764, 7765, 7764, 7764,
  5851, 5966, 5225, 5287, 5330, 5362, 5394, 5415, 5437, 5505, 5505, 5505, 
    5505, 5505, 5505, 6862, 7781, 7781, 7781, 7781, 7781, 7781,
  5211, 5498, 5542, 5580, 5607, 5627, 5647, 5660, 5675, 5718, 5718, 5718, 
    5718, 5718, 5718, 6884, 7281, 7436, 7436, 7436, 7436, 7436,
  4991, 5238, 5401, 5436, 5460, 5479, 5497, 5509, 5523, 5563, 5563, 5563, 
    5563, 5563, 5563, 6510, 7057, 7211, 7211, 7211, 7211, 7211,
  5096, 5370, 5476, 5513, 5539, 5559, 5578, 5591, 5606, 5648, 5648, 5648, 
    5648, 5648, 5648, 6718, 7189, 7343, 7343, 7343, 7343, 7343,
  5401, 5663, 5661, 5696, 5721, 5740, 5758, 5770, 5784, 5824, 5824, 5824, 
    5824, 5824, 5824, 6940, 7290, 7440, 7440, 7440, 7440, 7440,
  5765, 6015, 5962, 5994, 6017, 6035, 6051, 6063, 6075, 6112, 6112, 6112, 
    6112, 6112, 6112, 7202, 7470, 7612, 7612, 7612, 7612, 7612,
  6113, 6346, 6341, 6370, 6391, 6406, 6421, 6431, 6443, 6476, 6476, 6476, 
    6476, 6476, 6476, 7413, 7685, 7815, 7815, 7815, 7815, 7815,
  6409, 6646, 6752, 6779, 6799, 6814, 6829, 6838, 6849, 6881, 6881, 6881, 
    6881, 6881, 6881, 7667, 7988, 8108, 8108, 8108, 8108, 8108,
  6657, 6880, 6965, 6990, 7008, 7022, 7035, 7044, 7054, 7083, 7083, 7083, 
    7083, 7083, 7083, 7814, 8094, 8207, 8207, 8207, 8207, 8207,
  6756, 6986, 6970, 6996, 7015, 7029, 7043, 7051, 7062, 7091, 7091, 7091, 
    7091, 7091, 7091, 7946, 8124, 8238, 8238, 8238, 8238, 8238,
  6791, 7018, 6925, 6951, 6970, 6984, 6997, 7006, 7016, 7045, 7045, 7045, 
    7045, 7045, 7045, 7972, 8086, 8201, 8201, 8201, 8201, 8201,
  6671, 6879, 6687, 6712, 6730, 6743, 6756, 6765, 6775, 6803, 6803, 6803, 
    6803, 6803, 6803, 7809, 7872, 7993, 7993, 7993, 7993, 7993,
  6507, 6730, 6581, 6607, 6627, 6641, 6655, 6664, 6675, 6706, 6706, 6706, 
    6706, 6706, 6706, 7727, 7838, 7963, 7963, 7963, 7963, 7963,
  6286, 6512, 6397, 6425, 6445, 6460, 6474, 6484, 6495, 6527, 6527, 6527, 
    6527, 6527, 6527, 7548, 7714, 7844, 7844, 7844, 7844, 7844,
  6027, 6261, 6140, 6170, 6191, 6208, 6223, 6233, 6245, 6280, 6280, 6280, 
    6280, 6280, 6280, 7366, 7555, 7691, 7691, 7691, 7691, 7691,
  5814, 6071, 6011, 6044, 6067, 6085, 6102, 6113, 6126, 6163, 6163, 6163, 
    6163, 6163, 6163, 7270, 7520, 7661, 7661, 7661, 7661, 7661,
  5545, 5818, 5726, 5762, 5787, 5806, 5825, 5837, 5851, 5892, 5892, 5892, 
    5892, 5892, 5892, 7121, 7369, 7519, 7519, 7519, 7519, 7519,
  5251, 5529, 5439, 5476, 5502, 5523, 5542, 5555, 5569, 5613, 5613, 5613, 
    5613, 5613, 5613, 6895, 7181, 7339, 7339, 7339, 7339, 7339,
  5000, 5278, 5219, 5257, 5284, 5305, 5325, 5338, 5353, 5397, 5397, 5397, 
    5397, 5397, 5397, 6680, 7023, 7186, 7186, 7186, 7186, 7186,
  4895, 5184, 5168, 5208, 5236, 5257, 5278, 5292, 5307, 5353, 5353, 5353, 
    5353, 5353, 5353, 6632, 7018, 7182, 7182, 7182, 7182, 7182,
  5016, 5293, 5245, 5283, 5310, 5331, 5350, 5364, 5378, 5422, 5422, 5422, 
    5422, 5422, 5422, 6689, 7039, 7201, 7201, 7201, 7201, 7201,
  5360, 5637, 5612, 5648, 5674, 5694, 5713, 5726, 5740, 5782, 5782, 5782, 
    5782, 5782, 5782, 6976, 7299, 7452, 7452, 7452, 7452, 7452,
  5909, 6171, 6232, 6265, 6288, 6305, 6322, 6333, 6346, 6383, 6383, 6383, 
    6383, 6383, 6383, 7357, 7690, 7825, 7825, 7825, 7825, 7825,
  6528, 6746, 6912, 6937, 6955, 6969, 6982, 6991, 7001, 7030, 7030, 7030, 
    7030, 7030, 7030, 7675, 8042, 8155, 8155, 8155, 8155, 8155,
  7149, 7330, 7513, 7532, 7546, 7556, 7566, 7572, 7580, 7601, 7601, 7601, 
    7601, 7601, 7601, 8038, 8361, 8456, 8456, 8456, 8456, 8456,
  7690, 7967, 8056, 8065, 8072, 8077, 8081, 8084, 8087, 8098, 8098, 8098, 
    8098, 8098, 8098, 8492, 8439, 8439, 8439, 8439, 8440, 8439,
  7840, 8059, 8034, 8041, 8045, 8049, 8052, 8054, 8056, 8064, 8064, 8064, 
    8064, 8064, 8064, 8365, 8304, 8303, 8303, 8304, 8304, 8304,
  7981, 8177, 8114, 8118, 8121, 8123, 8125, 8126, 8128, 8132, 8132, 8132, 
    8132, 8132, 8132, 8375, 8277, 8277, 8277, 8277, 8277, 8277,
  7912, 8034, 8095, 8105, 8113, 8118, 8124, 8127, 8132, 8143, 8143, 8143, 
    8143, 8143, 8143, 8442, 8605, 8681, 8681, 8681, 8681, 8681,
  7735, 7902, 8176, 8186, 8193, 8198, 8204, 8207, 8210, 8221, 8221, 8221, 
    8221, 8221, 8221, 8429, 8590, 8590, 8590, 8590, 8590, 8590,
  7838, 8000, 8345, 8351, 8356, 8359, 8364, 8366, 8368, 8376, 8376, 8376, 
    8376, 8376, 8376, 8510, 8633, 8633, 8633, 8633, 8633, 8633,
  7866, 8299, 8728, 8721, 8716, 8711, 8707, 8704, 8701, 8693, 8693, 8693, 
    8693, 8693, 8693, 9026, 8403, 8403, 8403, 8403, 8403, 8403,
  7797, 7948, 8188, 8201, 8210, 8217, 8224, 8228, 8234, 8249, 8249, 8249, 
    8249, 8249, 8249, 8445, 8750, 8825, 8825, 8825, 8825, 8825,
  7330, 7581, 7867, 7862, 7858, 7855, 7852, 7850, 7848, 7841, 7841, 7841, 
    7841, 7841, 7841, 7763, 7631, 7631, 7631, 7631, 7631, 7631,
  6896, 7206, 7683, 7675, 7670, 7666, 7662, 7659, 7657, 7648, 7648, 7648, 
    7648, 7648, 7648, 7528, 7365, 7365, 7365, 7365, 7365, 7365,
  6917, 7124, 8014, 8034, 8049, 8060, 8070, 8077, 8085, 8107, 8107, 8107, 
    8107, 8107, 8107, 7851, 8765, 8842, 8842, 8842, 8842, 8842 ;

 Freq = 23.8, 31.4, 50.3, 51.76, 52.8, 53.596, 54.4, 54.94, 55.5, 57.29, 
    57.29, 57.29, 57.29, 57.29, 57.29, 88.2, 165.5, 183.31, 183.31, 183.31, 
    183.31, 183.31 ;

 GWP =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, _, _, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 0, 0, 0, 0, 0, 
    0, 24, 23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, _, _, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 20, 0, 0, 23, 24, 19, 21, 
    20, 0, 29, 44, 41, 33, 0, 35, 28, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, _, _, _, _, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, 
    _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 0, 0, 21, 0, 
    0, 0, 33, 35, 32, 30, 19, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, _, _, _, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 0, 0, 19, 24, 0, 0, 0, 21, 
    22, 0, 0, 0, 25, 24, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, _, _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 21, 25, 25, 23, 21, 23, 25, 26, 22, 0, 27, 24, 0, 0, 
    27, 32, 0, 26, 26, 25, 0, 17, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, _, _, 0, 0, 0, 0, _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 27, 31, 30, 25, 26, 24, 0, 0, 0, 25, 27, 29, 32, 29, 
    33, 37, 29, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, _, _, _, _, 0, 0, _, _, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 28, 26, 0, 0, 0, 0, 33, 38, 33, 34, 32, 
    29, 21, 21, 24, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 28, 33, 30, 27, 24, 
    23, 24, 21, 0, 0, 13, 0, 0, 0, 0, 0, 0, 0, 0, _, 0, 0, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 11, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 21, 0, 0, 0, 0, 0, 29, 26, 0, 
    22, 24, 22, 0, 0, 14, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 0, 0, 0, _, _, _, _, 
    _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 15, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 0, 0, 0, 0, 0, 0, 0, 0, 16, 17, 
    20, 22, 0, 0, 16, 15, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 0, 0, 0, _, _, _, 
    _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 16, 16, 10, 0, 12, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 
    21, 25, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 0, 0, _, _, _, _, _ ;

 IWP =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 LWP =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 
    1, 2, 1, 2, 2, 1, 1, 0, 2, 4, 6, 5, 24, 32, 60, 90, 60, 52, 58, 44, 42, 
    25, 27, 34, 46, 23, 27, 37, 70, 74, 83, 62, 31, 29, 5, 2, 1, 2, 1, 1, 3, 
    2, 1, 2, 1, 1, 4, 5, 10, 15, 0, -998, -998, 9, 13, 3, 1, 2, 6, 9, 14, 14, 
    2, -998, -998, -998, -998, -998, -998, -998, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 5, 5, 
    4, 3, 3, 7, 5, 6, 7, 15, 16, 25, 34, 44, 60, 71, 133, 172, 127, 38, 21, 
    109, 101, 132, 140, 129, 102, 22, 18, 87, 72, 98, 102, 37, 23, 8, 4, 2, 
    2, 2, 1, 2, 0, 1, 0, 0, 1, 1, 2, 4, 19, 8, 0, -998, -998, 2, 13, 6, 6, 
    11, 17, 24, 13, 4, -998, -998, -998, -998, -998, -998, -998, -998, -998,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 5, 7, 11, 
    7, 23, 9, 21, 33, 47, 56, 48, 45, 52, 47, 59, 58, 76, 20, 21, 75, 47, 17, 
    22, 18, 18, 19, 127, 16, 10, 13, 14, 138, 14, 11, 7, 0, 1, 2, 2, 2, 1, 1, 
    0, 1, 1, 1, 0, 1, 1, 3, 23, 17, -998, -998, -998, -998, 8, 12, 14, 18, 
    19, 19, 17, 9, -998, -998, -998, -998, -998, -998, -998, -998, -998, -998,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 2, 21, 18, 19, 
    8, 7, 28, 27, 32, 52, 48, 80, 58, 60, 54, 57, 41, 45, 59, 55, 52, 48, 34, 
    46, 14, 43, 53, 16, 43, 52, 83, 14, 13, 13, 10, 7, 6, 1, 0, 2, 2, 3, 1, 
    0, 0, 0, 0, 0, 2, 2, 4, 16, 16, 16, -998, -998, -998, 0, 10, 16, 21, 17, 
    14, 8, 7, -998, -998, -998, -998, -998, -998, -998, -998, -998, -998, -998,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 18, 26, 52, 36, 9, 4, 7, 
    10, 3, 4, 11, 19, 24, 29, 56, 52, 45, 50, 84, 98, 85, 72, 72, 20, 56, 52, 
    16, 18, 70, 54, 71, 13, 13, 43, 63, 73, 11, 8, 6, 28, 4, 3, 2, 1, 4, 3, 
    1, 1, 1, 0, 2, 2, 6, 12, 15, 13, 16, 16, 4, 1, -998, -998, 14, 20, 21, 
    -998, -998, -998, -998, -998, -998, -998, -998, -998, -998, -998, -998, 
    -998, -998, -998,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 3, 32, 80, 76, 44, 6, 4, 11, 
    10, 14, 15, 19, 33, 31, 30, 46, 54, 16, 18, 20, 21, 20, 19, 23, 18, 18, 
    55, 15, 10, 23, 70, 12, 12, 76, 9, 14, 10, 28, 6, 6, 8, 4, 3, 3, 2, 4, 2, 
    1, 0, 2, 2, 4, 8, 10, 17, 11, -998, -998, 9, 15, 15, 3, -998, 12, 16, 11, 
    -998, -998, -998, -998, -998, -998, -998, -998, -998, -998, -998, -998, 
    -998, -998, -998,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 29, 85, 63, 16, 12, 5, 3, 
    4, 12, 19, 30, 32, 24, 30, 51, 98, 15, 14, 17, 18, 17, 20, 135, 50, 41, 
    13, 14, 12, 11, 10, 9, 8, 10, 44, 66, 39, 31, 23, 5, 3, 1, 2, 3, 1, 4, 6, 
    9, 6, 8, 12, 13, 10, 10, 2, -998, -998, -998, -998, 17, 16, -998, -998, 
    0, -998, -998, -998, -998, -998, -998, -998, -998, -998, -998, -998, 
    -998, -998, -998, -998, -998, -998,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 7, 8, 24, 82, 26, 16, 13, 26, 20, 
    20, 21, 30, 50, 41, 31, 53, 63, 64, 92, 99, 87, 107, 16, 14, 73, 70, 78, 
    84, 12, 9, 10, 11, 10, 9, 8, 7, 8, 43, 27, 18, 4, 2, 1, 2, 2, 3, 3, 13, 
    11, 13, 13, 6, 11, 10, -998, -998, -998, -998, -998, -998, -998, -998, 
    -998, -998, -998, -998, -998, -998, -998, -998, -998, -998, -998, -998, 
    -998, -998, -998, -998, -998, -998, -998, -998,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 22, 37, 38, 26, 5, 3, 8, 16, 4, 
    20, 24, 24, 27, 35, 32, 44, 44, 43, 45, 45, 64, 55, 45, 60, 54, 46, 38, 
    58, 59, 11, 9, 8, 8, 7, 6, 6, 7, 27, 22, 4, 0, 0, 3, 3, 2, 7, 6, 6, -998, 
    11, 8, -998, -998, -998, -998, -998, -998, -998, -998, -998, -998, -998, 
    -998, -998, -998, -998, -998, -998, -998, -998, -998, -998, -998, -998, 
    0, 0, -998, -998, -998, -998, -998, -998,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 2, 20, 64, 12, 10, 38, 5, 4, 4, 7, 26, 
    16, 26, 26, 36, 26, 39, 34, 35, 30, 40, 44, 41, 49, 48, 8, 10, 43, 32, 
    27, 46, 72, 10, 9, 33, 7, 6, 8, 29, 23, 5, 1, 0, 1, 4, 8, 5, 8, 6, -998, 
    -998, -998, -998, -998, -998, -998, -998, -998, -998, -998, -998, -998, 
    -998, -998, -998, -998, -998, -998, -998, -998, -998, -998, -998, -998, 
    -998, 0, 0, 0, -998, -998, -998, -998, -998, -998,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 63, 37, 46, 14, 10, 44, 3, 2, 5, 36, 
    59, 40, 35, 34, 27, 37, 34, 15, 38, 40, 46, 44, 58, 52, 17, 54, 72, 59, 
    36, 22, 27, 23, 21, 5, 5, 6, 7, 24, 28, 7, 7, 4, 5, 4, 6, 9, 7, 5, -998, 
    -998, -998, -998, -998, -998, -998, -998, -998, -998, -998, -998, -998, 
    -998, -998, -998, -998, -998, -998, -998, -998, -998, -998, -998, -998, 
    -998, -998, -998, 0, 3, 6, -998, -998, -998, -998, -998,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 22, 9, 9, 9, 8, 101, 9, 36, 12, 3, 24, 38, 
    48, 42, 32, 33, 11, 28, 30, 38, 63, 40, 41, 67, 50, 61, 19, 44, 41, 54, 
    43, 31, 12, 13, 12, 2, 0, 6, 7, 6, 25, 17, 2, 8, 6, 4, 7, 8, 3, -998, 
    -998, -998, -998, -998, -998, -998, -998, -998, -998, -998, -998, -998, 
    -998, -998, -998, -998, -998, -998, -998, -998, -998, -998, -998, -998, 
    -998, -998, -998, -998, -998, 4, 7, -998, -998, -998, -998, -998 ;

 LZ_angle =
  -63.92, -62.21998, -60.58, -58.96998, -57.39001, -55.84999, -54.35999, 
    -52.89001, -51.41999, -49.96999, -48.53999, -47.15001, -45.77, -44.39001, 
    -42.98999, -41.60999, -40.27, -38.94, -37.60999, -36.28001, -34.95001, 
    -33.64001, -32.34001, -31.03001, -29.71, -28.41, -27.14001, -25.87, 
    -24.57999, -23.28, -22, -20.74, -19.48, -18.20999, -16.92, -15.65, -14.4, 
    -13.15, -11.88, -10.61, -9.36, -8.11, -6.86, -5.599999, -4.330001, 
    -3.080001, -1.85, -0.6000001, 0.6599999, 1.93, 3.19, 4.440001, 5.68, 
    6.940001, 8.22, 9.47, 10.72, 11.97, 13.25, 14.52, 15.78, 17.03, 18.3, 
    19.59, 20.87, 22.14001, 23.4, 24.67999, 25.98, 27.28, 28.57001, 29.85, 
    31.15, 32.46, 33.78001, 35.09001, 36.40999, 37.73999, 39.09001, 40.44, 
    41.78999, 43.14001, 44.51001, 45.91999, 47.33001, 48.73999, 50.15001, 
    51.58001, 53.07, 54.58001, 56.08001, 57.62, 59.18001, 60.81001, 62.47999, 
    64.18999,
  -63.96, -62.25, -60.59, -58.96998, -57.41, -55.90001, -54.39001, -52.90001, 
    -51.43, -49.98999, -48.57, -47.15999, -45.75, -44.34999, -42.98999, 
    -41.64001, -40.28999, -38.93, -37.59001, -36.28001, -34.96999, -33.65001, 
    -32.32, -31.01, -29.71, -28.44, -27.16, -25.85, -24.55, -23.28, -22.02, 
    -20.74, -19.47, -18.19, -16.92999, -15.68, -14.41, -13.13, -11.87, 
    -10.62, -9.380001, -8.119999, -6.839998, -5.580001, -4.339999, -3.099999, 
    -1.86, -0.58, 0.6800001, 1.93, 3.18, 4.440001, 5.699999, 6.960001, 
    8.199998, 9.449998, 10.72, 11.99, 13.26, 14.5, 15.76, 17.04001, 18.32001, 
    19.6, 20.85999, 22.12, 23.41, 24.7, 25.99, 27.26, 28.54999, 29.85, 31.16, 
    32.46, 33.76001, 35.07, 36.41999, 37.76001, 39.09999, 40.41999, 41.76001, 
    43.14001, 44.53999, 45.93, 47.31, 48.71999, 50.15001, 51.60999, 53.07, 
    54.55, 56.06001, 57.62, 59.21, 60.81001, 62.46, 64.16003,
  -63.96, -62.22999, -60.56999, -58.97999, -57.42, -55.88, -54.35999, -52.88, 
    -51.43, -50, -48.56, -47.14001, -45.73999, -44.37, -43.01001, -41.63, 
    -40.26001, -38.93, -37.60999, -36.29999, -34.96999, -33.63, -32.32, 
    -31.03001, -29.73, -28.42999, -27.13, -25.84, -24.57001, -23.3, -22.01, 
    -20.73, -19.45999, -18.20999, -16.95, -15.67, -14.39, -13.13, -11.89, 
    -10.64, -9.369999, -8.100001, -6.85, -5.599999, -4.36, -3.099999, -1.83, 
    -0.5900001, 0.6599999, 1.91, 3.19, 4.449999, 5.699999, 6.940001, 
    8.199998, 9.47, 10.74, 11.99, 13.24, 14.5, 15.77, 17.05, 18.31, 19.57001, 
    20.85, 22.14001, 23.42999, 24.69, 25.97, 27.26, 28.57001, 29.87, 31.15, 
    32.44, 33.76001, 35.09001, 36.41999, 37.75, 39.08001, 40.43, 41.79999, 
    43.16999, 44.53001, 45.90001, 47.31, 48.72999, 50.15999, 51.59001, 53.05, 
    54.55, 56.09, 57.64001, 59.18999, 60.79, 62.46998, 64.19999,
  -63.92, -62.21998, -60.59, -58.97999, -57.40001, -55.87, -54.37, -52.90001, 
    -51.43, -49.96999, -48.53999, -47.15001, -45.77, -44.38, -42.98999, 
    -41.60999, -40.28001, -38.95001, -37.62, -36.28001, -34.95001, -33.65001, 
    -32.34001, -31.03001, -29.71, -28.42, -27.14001, -25.87, -24.57001, 
    -23.28, -22, -20.74, -19.48, -18.2, -16.92999, -15.65, -14.4, -13.15, 
    -11.88, -10.62, -9.36, -8.119999, -6.87, -5.599999, -4.330001, -3.080001, 
    -1.84, -0.6000001, 0.67, 1.94, 3.19, 4.440001, 5.68, 6.949998, 8.22, 
    9.47, 10.73, 11.98, 13.25, 14.52, 15.78, 17.03, 18.29001, 19.57999, 
    20.87, 22.14001, 23.4, 24.67999, 25.97, 27.28, 28.57001, 29.85, 31.15, 
    32.46, 33.78001, 35.09001, 36.40001, 37.73999, 39.09999, 40.45001, 
    41.78999, 43.14001, 44.51001, 45.93, 47.33001, 48.73999, 50.15001, 
    51.59001, 53.07, 54.57, 56.08001, 57.59999, 59.18999, 60.81999, 62.47999, 
    64.18999,
  -63.96, -62.23999, -60.58, -58.96, -57.41, -55.89001, -54.39001, -52.89001, 
    -51.43, -49.98999, -48.57, -47.15999, -45.75, -44.35999, -43, -41.65001, 
    -40.28999, -38.93, -37.58001, -36.28001, -34.96999, -33.65001, -32.32, 
    -31, -29.71, -28.44, -27.15, -25.85, -24.55, -23.29001, -22.02, -20.74, 
    -19.47, -18.2, -16.94, -15.69, -14.41, -13.12, -11.86, -10.62, -9.369999, 
    -8.11, -6.839998, -5.580001, -4.349999, -3.11, -1.85, -0.58, 0.6800001, 
    1.92, 3.18, 4.440001, 5.71, 6.970001, 8.210002, 9.460003, 10.73, 12, 
    13.26, 14.5, 15.75, 17.03, 18.32001, 19.59, 20.85, 22.12, 23.41, 24.7, 
    25.99, 27.27, 28.56, 29.87, 31.17, 32.46999, 33.76001, 35.07, 36.41999, 
    37.77, 39.09999, 40.43, 41.77, 43.15001, 44.54999, 45.93, 47.31, 
    48.71999, 50.15001, 51.60999, 53.08001, 54.56001, 56.07, 57.64001, 
    59.21998, 60.81999, 62.45, 64.16003,
  -63.95, -62.21998, -60.56999, -58.98999, -57.43001, -55.89001, -54.37, 
    -52.89001, -51.43999, -50, -48.56, -47.13, -45.75, -44.38, -43.02, 
    -41.63, -40.26001, -38.93, -37.62, -36.29999, -34.96, -33.63, -32.32, 
    -31.03001, -29.73, -28.42999, -27.13, -25.85, -24.57001, -23.29001, -22, 
    -20.72, -19.47, -18.22, -16.95, -15.67, -14.39, -13.13, -11.89, -10.63, 
    -9.36, -8.089997, -6.85, -5.61, -4.36, -3.09, -1.83, -0.5900001, 
    0.6599999, 1.92, 3.2, 4.46, 5.699999, 6.940001, 8.199998, 9.479997, 
    10.74, 11.99, 13.24, 14.51, 15.78, 17.05, 18.3, 19.57001, 20.85, 
    22.14001, 23.42001, 24.69, 25.97, 27.26, 28.57001, 29.87, 31.15, 
    32.45001, 33.76001, 35.09999, 36.43, 37.73999, 39.07, 40.41999, 41.79999, 
    43.15999, 44.53001, 45.90001, 47.32, 48.75, 50.16999, 51.59001, 53.05, 
    54.56001, 56.09, 57.63, 59.18999, 60.79, 62.46998, 64.19999,
  -63.93001, -62.23999, -60.59, -58.97999, -57.40001, -55.87, -54.38, 
    -52.90001, -51.43, -49.96999, -48.53999, -47.15001, -45.77, -44.38, 
    -42.98999, -41.63, -40.28001, -38.95001, -37.60999, -36.27, -34.95001, 
    -33.65001, -32.34001, -31.02, -29.71, -28.42, -27.14001, -25.85999, 
    -24.57001, -23.27, -22, -20.74, -19.48, -18.2, -16.92, -15.67, -14.41, 
    -13.15, -11.88, -10.61, -9.350002, -8.119999, -6.86, -5.589998, 
    -4.330001, -3.09, -1.85, -0.6000001, 0.67, 1.94, 3.19, 4.43, 5.690001, 
    6.960001, 8.22, 9.47, 10.72, 11.98, 13.26, 14.52, 15.76, 17.02, 18.3, 
    19.59, 20.87, 22.14001, 23.4, 24.67999, 25.98, 27.28, 28.56, 29.85, 
    31.15, 32.46999, 33.78001, 35.09001, 36.40999, 37.75, 39.09999, 40.45001, 
    41.78999, 43.14001, 44.52, 45.91999, 47.33001, 48.72999, 50.15001, 
    51.59999, 53.08001, 54.58001, 56.08001, 57.60999, 59.18999, 60.81999, 
    62.47999, 64.17001,
  -63.96, -62.23999, -60.58, -58.97999, -57.42, -55.90001, -54.39001, 
    -52.89001, -51.41999, -49.98999, -48.57, -47.15001, -45.75, -44.35999, 
    -43, -41.65001, -40.28999, -38.91999, -37.59001, -36.28001, -34.96999, 
    -33.65001, -32.32, -31.01, -29.73, -28.44, -27.15, -25.84, -24.55, 
    -23.29001, -22.02, -20.74, -19.45999, -18.2, -16.94, -15.68, -14.4, 
    -13.12, -11.86, -10.62, -9.380001, -8.11, -6.839998, -5.589998, 
    -4.349999, -3.099999, -1.84, -0.58, 0.6800001, 1.92, 3.18, 4.440001, 
    5.71, 6.960001, 8.199998, 9.449998, 10.73, 12.01, 13.26, 14.51, 15.76, 
    17.04001, 18.32001, 19.59, 20.85, 22.12, 23.41, 24.7, 25.98, 27.26, 
    28.56, 29.87, 31.17, 32.46999, 33.76001, 35.08001, 36.41999, 37.77, 
    39.09001, 40.41999, 41.78001, 43.15999, 44.54999, 45.91999, 47.31, 
    48.71999, 50.16999, 51.62, 53.08001, 54.55, 56.08001, 57.64001, 59.21, 
    60.81001, 62.45, 64.17001,
  -63.96, -62.23999, -60.59, -59, -57.43999, -55.89001, -54.37, -52.90001, 
    -51.45, -50, -48.56, -47.13, -45.75, -44.38, -43.01001, -41.63, -40.27, 
    -38.93, -37.62, -36.29, -34.95001, -33.63, -32.32, -31.03001, -29.73, 
    -28.42, -27.12, -25.85, -24.57999, -23.29001, -22, -20.72, -19.47, 
    -18.22, -16.94, -15.66, -14.39, -13.14, -11.89, -10.63, -9.36, -8.100001, 
    -6.86, -5.61, -4.349999, -3.080001, -1.83, -0.5900001, 0.6499999, 1.92, 
    3.19, 4.449999, 5.690001, 6.940001, 8.210002, 9.479997, 10.73, 11.98, 
    13.24, 14.51, 15.78, 17.05, 18.3, 19.57001, 20.85999, 22.14001, 23.42001, 
    24.67999, 25.97, 27.27, 28.57001, 29.87, 31.15, 32.45001, 33.77, 
    35.10999, 36.43, 37.75, 39.08001, 40.44, 41.79999, 43.15001, 44.51001, 
    45.90999, 47.33001, 48.75, 50.15999, 51.59001, 53.05, 54.56001, 56.09, 
    57.63, 59.18999, 60.8, 62.47999, 64.19999,
  -63.93999, -62.23999, -60.58, -58.96998, -57.39001, -55.87, -54.38, 
    -52.89001, -51.43, -49.96999, -48.56, -47.15999, -45.77, -44.37, 
    -42.98999, -41.63, -40.28999, -38.94, -37.59999, -36.26001, -34.95001, 
    -33.65001, -32.34001, -31.01, -29.71, -28.42, -27.15, -25.85999, 
    -24.57001, -23.27, -22.01, -20.75, -19.48, -18.2, -16.92, -15.67, -14.41, 
    -13.15, -11.87, -10.61, -9.36, -8.119999, -6.86, -5.589998, -4.330001, 
    -3.09, -1.85, -0.6000001, 0.67, 1.94, 3.19, 4.43, 5.690001, 6.960001, 
    8.22, 9.460003, 10.72, 11.98, 13.26, 14.52, 15.76, 17.02, 18.31, 19.6, 
    20.87, 22.13, 23.4, 24.67999, 25.99, 27.28, 28.56, 29.85, 31.15, 
    32.46999, 33.78001, 35.08001, 36.40999, 37.76001, 39.10999, 40.45001, 
    41.78001, 43.14001, 44.53001, 45.93, 47.33001, 48.72999, 50.15001, 
    51.59999, 53.08001, 54.57, 56.07, 57.60999, 59.2, 60.83, 62.47999, 
    64.17001,
  -63.96998, -62.23999, -60.58, -58.96998, -57.42, -55.90001, -54.39001, 
    -52.89001, -51.43, -50, -48.58001, -47.15001, -45.73999, -44.37, 
    -43.01001, -41.65001, -40.28001, -38.93, -37.59999, -36.29, -34.96999, 
    -33.64001, -32.31, -31.01, -29.73, -28.45001, -27.14001, -25.84, -24.56, 
    -23.29001, -22.02, -20.74, -19.45999, -18.2, -16.95, -15.68, -14.39, 
    -13.12, -11.87, -10.63, -9.380001, -8.11, -6.839998, -5.589998, 
    -4.349999, -3.099999, -1.84, -0.58, 0.6800001, 1.92, 3.18, 4.449999, 
    5.699999, 6.940001, 8.190001, 9.460003, 10.74, 12.01, 13.26, 14.49, 
    15.76, 17.04001, 18.32001, 19.59, 20.85, 22.12, 23.42001, 24.7, 25.97, 
    27.26, 28.56, 29.87, 31.17, 32.45001, 33.75, 35.08001, 36.43, 37.77, 
    39.09001, 40.43, 41.78999, 43.16999, 44.53999, 45.90999, 47.29999, 
    48.72999, 50.16999, 51.62, 53.06001, 54.55, 56.08001, 57.64001, 59.21, 
    60.8, 62.45, 64.18002,
  -63.93999, -62.21998, -60.59, -58.98999, -57.42, -55.87, -54.37, -52.90001, 
    -51.43999, -49.98999, -48.54999, -47.14001, -45.77, -44.39001, -43, 
    -41.62, -40.26001, -38.94, -37.62, -36.28001, -34.95001, -33.63, 
    -32.33001, -31.03001, -29.73, -28.42, -27.13, -25.85999, -24.57001, 
    -23.29001, -22, -20.73, -19.48, -18.22, -16.92999, -15.65, -14.39, 
    -13.14, -11.9, -10.63, -9.36, -8.11, -6.86, -5.61, -4.339999, -3.080001, 
    -1.83, -0.6000001, 0.6599999, 1.93, 3.19, 4.440001, 5.68, 6.940001, 
    8.210002, 9.479997, 10.73, 11.98, 13.24, 14.51, 15.78, 17.04001, 18.3, 
    19.57001, 20.87, 22.15, 23.41, 24.67999, 25.97, 27.28, 28.57001, 
    29.85999, 31.14001, 32.45001, 33.77, 35.09001, 36.40999, 37.73999, 
    39.09001, 40.45001, 41.79999, 43.15001, 44.51001, 45.90999, 47.33001, 
    48.73999, 50.15999, 51.59001, 53.07, 54.57, 56.09, 57.62, 59.18001, 
    60.81001, 62.48999, 64.19999 ;

 Latitude =
  61.18, 61.58, 61.95, 62.28, 62.58, 62.86, 63.11, 63.34, 63.56, 63.77, 
    63.96, 64.14, 64.31, 64.47, 64.63, 64.78, 64.91, 65.04, 65.17, 65.29, 
    65.41, 65.52, 65.63, 65.73, 65.83, 65.93, 66.02, 66.11, 66.2, 66.28, 
    66.37, 66.45, 66.52, 66.6, 66.68, 66.75, 66.82, 66.89, 66.96, 67.03, 
    67.09, 67.16, 67.22, 67.28, 67.35, 67.41, 67.47, 67.52, 67.58, 67.64, 
    67.7, 67.75, 67.81, 67.87, 67.92, 67.98, 68.03, 68.08, 68.14, 68.19, 
    68.24, 68.29, 68.34, 68.4, 68.45, 68.5, 68.55, 68.6, 68.65, 68.7, 68.75, 
    68.79, 68.84, 68.89, 68.94, 68.99, 69.03, 69.08, 69.12, 69.17, 69.21, 
    69.25, 69.29, 69.33, 69.37, 69.4, 69.43, 69.46, 69.49, 69.5, 69.52, 
    69.52, 69.52, 69.5, 69.47, 69.42,
  61.28, 61.69, 62.06, 62.39, 62.69, 62.97, 63.22, 63.46, 63.69, 63.89, 
    64.08, 64.27, 64.44, 64.6, 64.76, 64.9, 65.04, 65.17, 65.3, 65.42, 65.54, 
    65.65, 65.76, 65.86, 65.96, 66.06, 66.15, 66.25, 66.33, 66.42, 66.5, 
    66.58, 66.66, 66.74, 66.82, 66.89, 66.96, 67.03, 67.1, 67.17, 67.23, 
    67.3, 67.36, 67.43, 67.49, 67.55, 67.61, 67.67, 67.73, 67.79, 67.84, 
    67.9, 67.96, 68.01, 68.07, 68.12, 68.18, 68.23, 68.28, 68.34, 68.39, 
    68.44, 68.49, 68.55, 68.6, 68.65, 68.7, 68.75, 68.8, 68.85, 68.9, 68.95, 
    68.99, 69.04, 69.09, 69.14, 69.18, 69.23, 69.28, 69.32, 69.36, 69.41, 
    69.45, 69.49, 69.52, 69.56, 69.59, 69.62, 69.64, 69.66, 69.67, 69.68, 
    69.67, 69.66, 69.62, 69.57,
  61.39, 61.81, 62.18, 62.51, 62.81, 63.09, 63.35, 63.59, 63.81, 64.01, 
    64.21, 64.39, 64.57, 64.73, 64.88, 65.03, 65.17, 65.31, 65.43, 65.55, 
    65.67, 65.78, 65.89, 66, 66.1, 66.2, 66.29, 66.38, 66.47, 66.56, 66.64, 
    66.72, 66.8, 66.88, 66.95, 67.03, 67.1, 67.17, 67.24, 67.31, 67.38, 
    67.44, 67.51, 67.57, 67.63, 67.69, 67.75, 67.81, 67.87, 67.93, 67.99, 
    68.05, 68.1, 68.16, 68.21, 68.27, 68.32, 68.38, 68.43, 68.48, 68.54, 
    68.59, 68.64, 68.69, 68.75, 68.8, 68.85, 68.9, 68.95, 69, 69.05, 69.1, 
    69.15, 69.19, 69.24, 69.29, 69.34, 69.38, 69.43, 69.47, 69.52, 69.56, 
    69.6, 69.64, 69.68, 69.71, 69.74, 69.77, 69.8, 69.82, 69.83, 69.83, 
    69.83, 69.81, 69.78, 69.72,
  61.51, 61.92, 62.29, 62.62, 62.93, 63.21, 63.47, 63.7, 63.93, 64.14, 64.34, 
    64.52, 64.69, 64.85, 65.01, 65.16, 65.3, 65.43, 65.56, 65.68, 65.8, 
    65.92, 66.02, 66.13, 66.23, 66.33, 66.42, 66.52, 66.61, 66.69, 66.78, 
    66.86, 66.94, 67.02, 67.09, 67.17, 67.24, 67.31, 67.38, 67.45, 67.52, 
    67.58, 67.65, 67.71, 67.77, 67.84, 67.9, 67.96, 68.02, 68.08, 68.13, 
    68.19, 68.25, 68.3, 68.36, 68.42, 68.47, 68.52, 68.58, 68.63, 68.69, 
    68.74, 68.79, 68.84, 68.9, 68.95, 69, 69.05, 69.1, 69.15, 69.2, 69.25, 
    69.3, 69.35, 69.4, 69.44, 69.49, 69.54, 69.58, 69.63, 69.67, 69.71, 
    69.76, 69.8, 69.83, 69.87, 69.9, 69.93, 69.95, 69.97, 69.98, 69.99, 
    69.98, 69.96, 69.93, 69.88,
  61.62, 62.03, 62.41, 62.74, 63.05, 63.33, 63.58, 63.83, 64.05, 64.26, 
    64.46, 64.64, 64.82, 64.98, 65.14, 65.28, 65.43, 65.56, 65.69, 65.82, 
    65.93, 66.05, 66.16, 66.27, 66.37, 66.46, 66.56, 66.65, 66.74, 66.83, 
    66.91, 67, 67.08, 67.15, 67.23, 67.31, 67.38, 67.45, 67.52, 67.59, 67.66, 
    67.72, 67.79, 67.85, 67.92, 67.98, 68.04, 68.1, 68.16, 68.22, 68.28, 
    68.34, 68.39, 68.45, 68.51, 68.56, 68.62, 68.67, 68.73, 68.78, 68.83, 
    68.89, 68.94, 68.99, 69.04, 69.1, 69.15, 69.2, 69.25, 69.3, 69.35, 69.4, 
    69.45, 69.5, 69.55, 69.6, 69.64, 69.69, 69.74, 69.78, 69.83, 69.87, 
    69.91, 69.95, 69.99, 70.02, 70.05, 70.08, 70.11, 70.13, 70.14, 70.14, 
    70.14, 70.12, 70.09, 70.03,
  61.73, 62.15, 62.52, 62.85, 63.16, 63.44, 63.71, 63.95, 64.17, 64.38, 
    64.58, 64.77, 64.94, 65.11, 65.26, 65.41, 65.56, 65.69, 65.82, 65.94, 
    66.06, 66.18, 66.29, 66.4, 66.5, 66.6, 66.69, 66.79, 66.88, 66.96, 67.05, 
    67.13, 67.21, 67.29, 67.37, 67.44, 67.52, 67.59, 67.66, 67.73, 67.8, 
    67.87, 67.93, 67.99, 68.06, 68.12, 68.18, 68.24, 68.3, 68.36, 68.42, 
    68.48, 68.54, 68.6, 68.65, 68.71, 68.76, 68.82, 68.87, 68.93, 68.98, 
    69.04, 69.09, 69.14, 69.19, 69.25, 69.3, 69.35, 69.4, 69.45, 69.5, 69.55, 
    69.6, 69.65, 69.7, 69.75, 69.8, 69.84, 69.89, 69.94, 69.98, 70.02, 70.07, 
    70.11, 70.14, 70.18, 70.21, 70.24, 70.26, 70.28, 70.29, 70.3, 70.29, 
    70.27, 70.24, 70.18,
  61.84, 62.26, 62.63, 62.97, 63.28, 63.56, 63.82, 64.06, 64.29, 64.51, 
    64.71, 64.89, 65.06, 65.23, 65.39, 65.54, 65.68, 65.82, 65.95, 66.08, 
    66.2, 66.31, 66.42, 66.53, 66.63, 66.73, 66.83, 66.92, 67.01, 67.1, 
    67.19, 67.27, 67.35, 67.43, 67.51, 67.58, 67.66, 67.73, 67.8, 67.87, 
    67.94, 68.01, 68.07, 68.14, 68.2, 68.26, 68.32, 68.39, 68.45, 68.51, 
    68.57, 68.63, 68.68, 68.74, 68.8, 68.85, 68.91, 68.97, 69.02, 69.08, 
    69.13, 69.18, 69.24, 69.29, 69.34, 69.4, 69.45, 69.5, 69.55, 69.6, 69.65, 
    69.7, 69.75, 69.8, 69.85, 69.9, 69.95, 70, 70.05, 70.09, 70.14, 70.18, 
    70.22, 70.26, 70.3, 70.33, 70.37, 70.39, 70.42, 70.44, 70.45, 70.45, 
    70.45, 70.43, 70.39, 70.34,
  61.94, 62.37, 62.74, 63.08, 63.39, 63.67, 63.94, 64.19, 64.41, 64.63, 
    64.82, 65.01, 65.19, 65.36, 65.52, 65.67, 65.81, 65.95, 66.08, 66.2, 
    66.32, 66.44, 66.55, 66.66, 66.76, 66.86, 66.96, 67.06, 67.15, 67.24, 
    67.32, 67.41, 67.49, 67.57, 67.64, 67.72, 67.8, 67.87, 67.94, 68.01, 
    68.08, 68.15, 68.21, 68.28, 68.34, 68.41, 68.47, 68.53, 68.59, 68.65, 
    68.71, 68.77, 68.83, 68.89, 68.94, 69, 69.06, 69.11, 69.17, 69.22, 69.28, 
    69.33, 69.39, 69.44, 69.49, 69.55, 69.6, 69.65, 69.7, 69.75, 69.81, 
    69.86, 69.91, 69.96, 70.01, 70.05, 70.1, 70.15, 70.2, 70.24, 70.29, 
    70.33, 70.38, 70.42, 70.45, 70.49, 70.52, 70.55, 70.57, 70.59, 70.6, 
    70.61, 70.6, 70.58, 70.55, 70.49,
  62.05, 62.48, 62.85, 63.19, 63.5, 63.79, 64.06, 64.3, 64.53, 64.74, 64.95, 
    65.14, 65.31, 65.48, 65.64, 65.79, 65.94, 66.08, 66.21, 66.33, 66.46, 
    66.57, 66.68, 66.79, 66.9, 67, 67.1, 67.19, 67.28, 67.37, 67.46, 67.54, 
    67.62, 67.7, 67.78, 67.86, 67.94, 68.01, 68.08, 68.15, 68.22, 68.29, 
    68.35, 68.42, 68.48, 68.55, 68.61, 68.67, 68.73, 68.8, 68.86, 68.92, 
    68.97, 69.03, 69.09, 69.15, 69.2, 69.26, 69.31, 69.37, 69.43, 69.48, 
    69.53, 69.59, 69.64, 69.7, 69.75, 69.8, 69.85, 69.9, 69.96, 70.01, 70.06, 
    70.11, 70.16, 70.21, 70.26, 70.3, 70.35, 70.4, 70.44, 70.49, 70.53, 
    70.57, 70.61, 70.64, 70.68, 70.7, 70.73, 70.75, 70.76, 70.76, 70.76, 
    70.74, 70.7, 70.64,
  62.17, 62.59, 62.97, 63.31, 63.63, 63.91, 64.18, 64.42, 64.65, 64.87, 
    65.07, 65.26, 65.44, 65.61, 65.77, 65.92, 66.06, 66.2, 66.34, 66.46, 
    66.58, 66.7, 66.81, 66.92, 67.03, 67.13, 67.23, 67.32, 67.42, 67.51, 
    67.59, 67.68, 67.76, 67.84, 67.92, 68, 68.07, 68.15, 68.22, 68.29, 68.36, 
    68.43, 68.49, 68.56, 68.63, 68.69, 68.75, 68.82, 68.88, 68.94, 69, 69.06, 
    69.12, 69.18, 69.24, 69.29, 69.35, 69.41, 69.46, 69.52, 69.57, 69.63, 
    69.68, 69.74, 69.79, 69.84, 69.9, 69.95, 70, 70.06, 70.11, 70.16, 70.21, 
    70.26, 70.31, 70.36, 70.41, 70.46, 70.51, 70.55, 70.6, 70.64, 70.68, 
    70.73, 70.76, 70.8, 70.83, 70.86, 70.88, 70.9, 70.91, 70.92, 70.91, 
    70.89, 70.85, 70.8,
  62.27, 62.7, 63.08, 63.43, 63.74, 64.02, 64.29, 64.54, 64.77, 64.99, 65.19, 
    65.38, 65.56, 65.73, 65.89, 66.04, 66.19, 66.33, 66.46, 66.59, 66.71, 
    66.83, 66.95, 67.06, 67.16, 67.26, 67.36, 67.46, 67.55, 67.64, 67.73, 
    67.81, 67.9, 67.98, 68.06, 68.13, 68.21, 68.29, 68.36, 68.43, 68.5, 
    68.57, 68.64, 68.7, 68.77, 68.83, 68.9, 68.96, 69.02, 69.08, 69.14, 69.2, 
    69.26, 69.32, 69.38, 69.44, 69.5, 69.55, 69.61, 69.66, 69.72, 69.78, 
    69.83, 69.89, 69.94, 69.99, 70.05, 70.1, 70.15, 70.21, 70.26, 70.31, 
    70.36, 70.41, 70.46, 70.51, 70.56, 70.61, 70.66, 70.71, 70.75, 70.8, 
    70.84, 70.88, 70.92, 70.95, 70.99, 71.02, 71.04, 71.06, 71.07, 71.07, 
    71.07, 71.05, 71.01, 70.95,
  62.38, 62.81, 63.19, 63.54, 63.85, 64.14, 64.41, 64.66, 64.89, 65.11, 
    65.31, 65.5, 65.68, 65.85, 66.02, 66.17, 66.32, 66.46, 66.59, 66.72, 
    66.84, 66.96, 67.08, 67.18, 67.29, 67.39, 67.49, 67.59, 67.68, 67.77, 
    67.86, 67.95, 68.03, 68.11, 68.19, 68.27, 68.35, 68.42, 68.5, 68.57, 
    68.64, 68.71, 68.77, 68.84, 68.91, 68.97, 69.04, 69.1, 69.16, 69.23, 
    69.29, 69.35, 69.41, 69.47, 69.53, 69.58, 69.64, 69.7, 69.75, 69.81, 
    69.87, 69.92, 69.98, 70.03, 70.09, 70.14, 70.2, 70.25, 70.3, 70.36, 
    70.41, 70.46, 70.51, 70.56, 70.62, 70.67, 70.72, 70.76, 70.81, 70.86, 
    70.91, 70.95, 70.99, 71.03, 71.07, 71.11, 71.14, 71.17, 71.2, 71.21, 
    71.23, 71.23, 71.22, 71.2, 71.16, 71.1 ;

 Longitude =
  135.75, 136.65, 137.5, 138.3, 139.06, 139.78, 140.45, 141.09, 141.71, 
    142.31, 142.89, 143.44, 143.97, 144.48, 144.99, 145.49, 145.96, 146.41, 
    146.86, 147.3, 147.73, 148.15, 148.56, 148.97, 149.37, 149.76, 150.14, 
    150.52, 150.9, 151.27, 151.64, 152, 152.35, 152.71, 153.07, 153.42, 
    153.77, 154.11, 154.46, 154.81, 155.15, 155.49, 155.83, 156.18, 156.53, 
    156.87, 157.21, 157.55, 157.9, 158.26, 158.61, 158.97, 159.32, 159.68, 
    160.05, 160.42, 160.79, 161.16, 161.55, 161.94, 162.33, 162.73, 163.14, 
    163.56, 163.99, 164.42, 164.85, 165.3, 165.77, 166.25, 166.73, 167.22, 
    167.74, 168.27, 168.82, 169.38, 169.96, 170.57, 171.2, 171.86, 172.53, 
    173.24, 173.98, 174.77, 175.59, 176.45, 177.34, 178.29, 179.32, -179.58, 
    -178.43, -177.2, -175.88, -174.42, -172.85, -171.14,
  135.49, 136.41, 137.26, 138.07, 138.82, 139.53, 140.2, 140.86, 141.49, 
    142.08, 142.65, 143.21, 143.75, 144.27, 144.77, 145.26, 145.73, 146.2, 
    146.65, 147.09, 147.51, 147.93, 148.35, 148.76, 149.16, 149.55, 149.93, 
    150.32, 150.7, 151.07, 151.43, 151.8, 152.16, 152.52, 152.87, 153.22, 
    153.57, 153.93, 154.27, 154.62, 154.96, 155.3, 155.65, 156, 156.34, 
    156.68, 157.03, 157.38, 157.74, 158.09, 158.44, 158.8, 159.16, 159.52, 
    159.89, 160.25, 160.63, 161.01, 161.4, 161.78, 162.18, 162.58, 163, 
    163.42, 163.84, 164.27, 164.72, 165.18, 165.64, 166.11, 166.6, 167.1, 
    167.63, 168.16, 168.7, 169.27, 169.86, 170.48, 171.11, 171.76, 172.44, 
    173.16, 173.92, 174.71, 175.52, 176.38, 177.29, 178.27, 179.29, -179.63, 
    -178.47, -177.21, -175.86, -174.41, -172.85, -171.13,
  135.26, 136.19, 137.04, 137.83, 138.58, 139.3, 139.99, 140.64, 141.25, 
    141.85, 142.43, 142.99, 143.53, 144.04, 144.54, 145.03, 145.52, 145.98, 
    146.42, 146.86, 147.3, 147.72, 148.14, 148.54, 148.94, 149.34, 149.73, 
    150.11, 150.49, 150.86, 151.23, 151.6, 151.96, 152.31, 152.67, 153.03, 
    153.38, 153.73, 154.07, 154.42, 154.77, 155.12, 155.47, 155.81, 156.16, 
    156.5, 156.86, 157.2, 157.55, 157.91, 158.27, 158.63, 158.99, 159.35, 
    159.72, 160.1, 160.48, 160.85, 161.24, 161.63, 162.03, 162.44, 162.85, 
    163.26, 163.69, 164.14, 164.59, 165.04, 165.5, 165.98, 166.48, 166.99, 
    167.5, 168.04, 168.59, 169.17, 169.76, 170.38, 171.01, 171.67, 172.37, 
    173.1, 173.84, 174.62, 175.45, 176.33, 177.25, 178.21, 179.24, -179.66, 
    -178.47, -177.2, -175.87, -174.42, -172.82, -171.06,
  135.04, 135.95, 136.8, 137.6, 138.36, 139.07, 139.75, 140.4, 141.02, 
    141.63, 142.21, 142.76, 143.29, 143.81, 144.32, 144.82, 145.29, 145.75, 
    146.2, 146.65, 147.08, 147.5, 147.92, 148.33, 148.74, 149.13, 149.52, 
    149.9, 150.28, 150.66, 151.03, 151.39, 151.75, 152.11, 152.47, 152.83, 
    153.18, 153.53, 153.88, 154.23, 154.58, 154.93, 155.27, 155.62, 155.98, 
    156.33, 156.67, 157.02, 157.38, 157.74, 158.1, 158.45, 158.81, 159.18, 
    159.56, 159.93, 160.31, 160.69, 161.08, 161.48, 161.88, 162.28, 162.69, 
    163.12, 163.56, 164, 164.44, 164.9, 165.37, 165.86, 166.36, 166.86, 
    167.38, 167.93, 168.49, 169.06, 169.65, 170.27, 170.92, 171.59, 172.28, 
    173, 173.75, 174.56, 175.4, 176.28, 177.19, 178.16, 179.21, -179.67, 
    -178.5, -177.24, -175.88, -174.39, -172.78, -171.03,
  134.79, 135.71, 136.56, 137.37, 138.12, 138.83, 139.51, 140.16, 140.79, 
    141.39, 141.96, 142.52, 143.07, 143.59, 144.09, 144.58, 145.06, 145.53, 
    145.99, 146.43, 146.85, 147.28, 147.71, 148.12, 148.52, 148.91, 149.3, 
    149.69, 150.07, 150.44, 150.81, 151.18, 151.55, 151.91, 152.27, 152.62, 
    152.98, 153.34, 153.69, 154.04, 154.38, 154.74, 155.09, 155.44, 155.79, 
    156.13, 156.49, 156.84, 157.2, 157.55, 157.91, 158.28, 158.65, 159.02, 
    159.39, 159.76, 160.14, 160.53, 160.92, 161.31, 161.71, 162.13, 162.55, 
    162.98, 163.41, 163.85, 164.3, 164.77, 165.24, 165.73, 166.22, 166.74, 
    167.27, 167.81, 168.36, 168.94, 169.55, 170.18, 170.83, 171.49, 172.19, 
    172.92, 173.7, 174.49, 175.33, 176.21, 177.14, 178.13, 179.18, -179.71, 
    -178.52, -177.23, -175.85, -174.37, -172.79, -171.02,
  134.56, 135.48, 136.33, 137.12, 137.87, 138.59, 139.28, 139.93, 140.55, 
    141.15, 141.74, 142.3, 142.83, 143.35, 143.85, 144.35, 144.84, 145.3, 
    145.75, 146.19, 146.63, 147.07, 147.49, 147.89, 148.29, 148.7, 149.09, 
    149.47, 149.85, 150.23, 150.61, 150.98, 151.34, 151.7, 152.06, 152.42, 
    152.78, 153.14, 153.48, 153.84, 154.19, 154.55, 154.89, 155.24, 155.59, 
    155.95, 156.31, 156.66, 157.01, 157.37, 157.74, 158.11, 158.47, 158.84, 
    159.21, 159.6, 159.98, 160.37, 160.76, 161.16, 161.56, 161.98, 162.39, 
    162.82, 163.26, 163.71, 164.16, 164.63, 165.1, 165.59, 166.1, 166.62, 
    167.14, 167.68, 168.25, 168.84, 169.45, 170.07, 170.72, 171.4, 172.11, 
    172.85, 173.61, 174.41, 175.26, 176.16, 177.1, 178.08, 179.13, -179.74, 
    -178.52, -177.24, -175.87, -174.39, -172.75, -170.95,
  134.33, 135.23, 136.08, 136.88, 137.64, 138.36, 139.04, 139.69, 140.32, 
    140.93, 141.51, 142.06, 142.59, 143.12, 143.63, 144.13, 144.6, 145.07, 
    145.53, 145.98, 146.41, 146.83, 147.25, 147.67, 148.08, 148.48, 148.87, 
    149.25, 149.64, 150.02, 150.39, 150.76, 151.13, 151.49, 151.86, 152.22, 
    152.57, 152.93, 153.29, 153.64, 154, 154.34, 154.7, 155.05, 155.41, 
    155.76, 156.11, 156.47, 156.83, 157.2, 157.56, 157.92, 158.29, 158.67, 
    159.05, 159.42, 159.81, 160.2, 160.6, 161, 161.4, 161.81, 162.24, 162.68, 
    163.12, 163.56, 164.01, 164.48, 164.97, 165.46, 165.96, 166.48, 167.01, 
    167.57, 168.14, 168.73, 169.33, 169.97, 170.63, 171.31, 172.02, 172.75, 
    173.53, 174.35, 175.2, 176.09, 177.04, 178.04, 179.12, -179.75, -178.55, 
    -177.26, -175.87, -174.35, -172.71, -170.94,
  134.07, 134.98, 135.84, 136.64, 137.39, 138.1, 138.79, 139.45, 140.08, 
    140.68, 141.26, 141.82, 142.36, 142.89, 143.39, 143.88, 144.37, 144.84, 
    145.3, 145.74, 146.18, 146.61, 147.04, 147.45, 147.85, 148.25, 148.65, 
    149.04, 149.43, 149.8, 150.18, 150.55, 150.92, 151.28, 151.64, 152, 
    152.37, 152.73, 153.09, 153.44, 153.79, 154.15, 154.5, 154.86, 155.21, 
    155.56, 155.93, 156.29, 156.65, 157.01, 157.37, 157.74, 158.12, 158.49, 
    158.86, 159.24, 159.64, 160.04, 160.43, 160.83, 161.24, 161.66, 162.09, 
    162.52, 162.96, 163.41, 163.87, 164.35, 164.83, 165.32, 165.83, 166.36, 
    166.9, 167.45, 168.01, 168.61, 169.23, 169.87, 170.53, 171.2, 171.92, 
    172.68, 173.46, 174.27, 175.12, 176.03, 177, 178.01, 179.07, -179.8, 
    -178.57, -177.25, -175.85, -174.34, -172.71, -170.9,
  133.83, 134.74, 135.59, 136.38, 137.14, 137.87, 138.55, 139.21, 139.83, 
    140.43, 141.02, 141.59, 142.12, 142.64, 143.15, 143.65, 144.14, 144.61, 
    145.06, 145.51, 145.95, 146.39, 146.81, 147.22, 147.62, 148.03, 148.43, 
    148.82, 149.2, 149.58, 149.96, 150.34, 150.7, 151.06, 151.43, 151.8, 
    152.16, 152.52, 152.87, 153.23, 153.59, 153.95, 154.3, 154.65, 155.01, 
    155.38, 155.73, 156.09, 156.45, 156.82, 157.19, 157.56, 157.93, 158.31, 
    158.69, 159.08, 159.47, 159.86, 160.26, 160.66, 161.08, 161.5, 161.92, 
    162.36, 162.81, 163.27, 163.73, 164.2, 164.68, 165.19, 165.7, 166.23, 
    166.76, 167.32, 167.9, 168.51, 169.12, 169.76, 170.42, 171.12, 171.84, 
    172.59, 173.36, 174.19, 175.07, 175.99, 176.94, 177.94, 179.02, -179.81, 
    -178.57, -177.27, -175.86, -174.33, -172.66, -170.83,
  133.59, 134.5, 135.35, 136.15, 136.92, 137.63, 138.31, 138.96, 139.59, 
    140.2, 140.78, 141.33, 141.88, 142.41, 142.92, 143.42, 143.9, 144.37, 
    144.83, 145.28, 145.72, 146.15, 146.57, 146.99, 147.41, 147.81, 148.2, 
    148.59, 148.98, 149.37, 149.74, 150.11, 150.48, 150.85, 151.22, 151.58, 
    151.95, 152.31, 152.67, 153.03, 153.39, 153.74, 154.1, 154.46, 154.82, 
    155.18, 155.53, 155.9, 156.26, 156.63, 157, 157.37, 157.75, 158.13, 
    158.51, 158.9, 159.29, 159.69, 160.09, 160.5, 160.91, 161.33, 161.76, 
    162.21, 162.66, 163.11, 163.57, 164.05, 164.55, 165.05, 165.56, 166.09, 
    166.64, 167.2, 167.78, 168.38, 169, 169.65, 170.33, 171.02, 171.74, 
    172.49, 173.29, 174.13, 175.01, 175.91, 176.88, 177.91, 179, -179.84, 
    -178.61, -177.29, -175.85, -174.3, -172.63, -170.82,
  133.33, 134.25, 135.11, 135.91, 136.66, 137.37, 138.06, 138.72, 139.35, 
    139.95, 140.53, 141.09, 141.64, 142.17, 142.67, 143.17, 143.66, 144.14, 
    144.59, 145.04, 145.48, 145.92, 146.35, 146.76, 147.17, 147.57, 147.97, 
    148.37, 148.76, 149.14, 149.52, 149.89, 150.27, 150.63, 151, 151.37, 
    151.74, 152.1, 152.46, 152.81, 153.17, 153.54, 153.9, 154.26, 154.61, 
    154.97, 155.34, 155.71, 156.07, 156.44, 156.81, 157.19, 157.57, 157.94, 
    158.32, 158.71, 159.12, 159.52, 159.92, 160.32, 160.74, 161.17, 161.61, 
    162.05, 162.49, 162.95, 163.43, 163.91, 164.4, 164.9, 165.42, 165.96, 
    166.51, 167.07, 167.65, 168.26, 168.9, 169.55, 170.22, 170.91, 171.65, 
    172.42, 173.22, 174.05, 174.92, 175.85, 176.84, 177.87, 178.95, -179.88, 
    -178.62, -177.27, -175.84, -174.3, -172.63, -170.76,
  133.09, 134.01, 134.85, 135.65, 136.41, 137.13, 137.81, 138.47, 139.09, 
    139.7, 140.29, 140.85, 141.39, 141.91, 142.43, 142.94, 143.42, 143.89, 
    144.35, 144.8, 145.25, 145.68, 146.11, 146.52, 146.94, 147.35, 147.74, 
    148.13, 148.52, 148.91, 149.3, 149.67, 150.04, 150.41, 150.78, 151.16, 
    151.52, 151.88, 152.24, 152.6, 152.97, 153.33, 153.69, 154.05, 154.41, 
    154.78, 155.14, 155.5, 155.87, 156.24, 156.62, 157, 157.37, 157.75, 
    158.14, 158.54, 158.93, 159.33, 159.74, 160.16, 160.58, 161, 161.43, 
    161.88, 162.34, 162.8, 163.27, 163.75, 164.25, 164.76, 165.29, 165.82, 
    166.37, 166.94, 167.53, 168.14, 168.77, 169.43, 170.11, 170.82, 171.56, 
    172.32, 173.12, 173.97, 174.86, 175.8, 176.78, 177.81, 178.92, -179.89, 
    -178.63, -177.3, -175.86, -174.28, -172.56, -170.7 ;

 Orb_mode = 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 Polo = 2, 2, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 2, 3, 3, 3, 3, 3, 3 ;

 PrecipType =
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888 ;

 Prob_SF =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, _, _, _, _, 0, 0, 0, 0, 0, 0, 0, 22, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 54, _, _, _, _, 0, 0, 0, 0, 0, 0, 10, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, _, _, _, _, _, _, 0, 0, 0, 16, 12, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    _, _, _, _, _, _, 0, 0, 20, 28, 48, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 27, 40, 
    _, _, _, _, _, 8, 0, 12, 33, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 28, 26, _, 
    _, 22, _, _, _, _, 12, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 30, _, _, _, _, 
    _, _, 23, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 65, 65, 0, 65, 65, 0, _, 63, 62, 51, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 65, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 65, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 64, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 39, _, _, _, _, _, _ ;

 Qc =
  1, 0, 144, 8192,
  1, 0, 144, 8192,
  1, 0, 144, 8192,
  1, 0, 144, 8192,
  0, 0, 128, 8192,
  1, 0, 144, 8192,
  0, 0, 128, 8192,
  0, 0, 128, 8192,
  1, 0, 144, 8192,
  1, 0, 144, 8192,
  1, 0, 144, 8192,
  0, 0, 128, 8192,
  0, 0, 128, 8192,
  0, 0, 128, 8192,
  1, 0, 156, 8192,
  0, 0, 128, 8192,
  0, 0, 128, 8192,
  0, 0, 128, 8192,
  0, 0, 128, 8192,
  0, 0, 128, 8192,
  0, 0, 128, 8192,
  0, 0, 128, 8192,
  0, 0, 128, 8192,
  0, 0, 160, 8192,
  0, 0, 160, 8192,
  0, 0, 128, 8192,
  0, 0, 160, 8192,
  1, 0, 148, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 148, 8192,
  1, 0, 140, 8192,
  1, 0, 156, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 180, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  0, 0, 160, 8192,
  1, 0, 180, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  0, 0, 160, 8192,
  1, 0, 164, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 180, 8192,
  1, 0, 176, 8192,
  1, 0, 176, 8192,
  1, 0, 176, 8192,
  1, 0, 188, 8192,
  1, 0, 172, 8192,
  0, 0, 128, 8192,
  0, 0, 160, 8192,
  0, 0, 128, 8192,
  0, 0, 128, 8192,
  0, 0, 160, 8192,
  0, 0, 160, 8192,
  0, 0, 128, 8192,
  0, 0, 160, 8192,
  0, 0, 128, 8192,
  0, 0, 128, 8192,
  0, 0, 160, 8192,
  0, 0, 160, 8192,
  0, 0, 160, 8192,
  0, 0, 160, 8192,
  1, 0, 144, 8192,
  0, 0, 128, 0,
  0, 0, 128, 0,
  1, 0, 176, 8192,
  0, 0, 160, 8192,
  0, 0, 160, 8192,
  0, 0, 128, 8192,
  0, 0, 160, 8192,
  0, 0, 160, 8192,
  0, 0, 160, 8192,
  0, 0, 160, 8192,
  0, 0, 160, 8192,
  0, 0, 160, 8192,
  0, 0, 128, 0,
  0, 0, 128, 0,
  0, 0, 128, 0,
  0, 0, 0, 4096,
  0, 0, 32, 4096,
  0, 0, 32, 4096,
  0, 0, 0, 4096,
  0, 0, 128, 0,
  1, 0, 144, 8192,
  1, 0, 144, 8192,
  0, 0, 128, 8192,
  1, 0, 144, 8192,
  1, 0, 144, 8192,
  1, 0, 144, 8192,
  1, 0, 144, 8192,
  1, 0, 148, 8192,
  0, 0, 128, 8192,
  1, 0, 144, 8192,
  1, 0, 144, 8192,
  0, 0, 128, 8192,
  0, 0, 128, 8192,
  1, 0, 144, 8192,
  0, 0, 128, 8192,
  0, 0, 128, 8192,
  0, 0, 128, 8192,
  0, 0, 128, 8192,
  0, 0, 128, 8192,
  0, 0, 128, 8192,
  0, 0, 128, 8192,
  0, 0, 128, 8192,
  0, 0, 160, 8192,
  0, 0, 160, 8192,
  1, 0, 180, 8192,
  0, 0, 160, 8192,
  0, 0, 160, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 172, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  0, 0, 160, 8192,
  1, 28, 3776, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 28, 3776, 8192,
  1, 12, 3776, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  0, 0, 160, 8192,
  1, 0, 176, 8192,
  1, 0, 188, 8192,
  1, 0, 180, 8192,
  0, 0, 160, 8192,
  0, 0, 160, 8192,
  0, 0, 160, 8192,
  0, 0, 128, 8192,
  0, 0, 160, 8192,
  0, 0, 128, 8192,
  0, 0, 128, 8192,
  0, 0, 128, 8192,
  0, 0, 128, 8192,
  0, 0, 128, 8192,
  0, 0, 128, 8192,
  0, 0, 160, 8192,
  0, 0, 160, 8192,
  1, 0, 176, 8192,
  1, 0, 176, 8192,
  1, 0, 144, 8192,
  0, 0, 128, 0,
  0, 0, 128, 0,
  0, 0, 160, 8192,
  0, 0, 160, 8192,
  0, 0, 160, 8192,
  0, 0, 160, 8192,
  0, 0, 160, 8192,
  0, 0, 160, 8192,
  0, 0, 160, 8192,
  0, 0, 160, 8192,
  0, 0, 160, 8192,
  0, 0, 128, 0,
  0, 0, 128, 0,
  0, 0, 128, 0,
  0, 0, 128, 0,
  0, 0, 0, 4096,
  0, 0, 32, 4096,
  0, 0, 0, 4096,
  0, 0, 0, 4096,
  1, 0, 28, 4096,
  1, 0, 144, 8192,
  1, 0, 144, 8192,
  1, 0, 144, 8192,
  1, 0, 144, 8192,
  1, 0, 144, 8192,
  1, 0, 144, 8192,
  1, 0, 144, 8192,
  1, 0, 144, 8192,
  1, 0, 144, 8192,
  1, 0, 148, 8192,
  1, 0, 144, 8192,
  1, 0, 148, 8192,
  1, 0, 144, 8192,
  1, 0, 144, 8192,
  0, 0, 128, 8192,
  0, 0, 128, 8192,
  0, 0, 128, 8192,
  0, 0, 128, 8192,
  0, 0, 128, 8192,
  0, 0, 128, 8192,
  0, 0, 128, 8192,
  0, 0, 160, 8192,
  1, 0, 164, 8192,
  1, 0, 180, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  0, 0, 160, 8192,
  1, 0, 188, 8192,
  1, 0, 164, 8192,
  1, 0, 180, 8192,
  1, 0, 180, 8192,
  1, 0, 180, 8192,
  1, 28, 3776, 8192,
  1, 28, 3776, 8192,
  1, 0, 180, 8192,
  0, 0, 160, 8192,
  1, 12, 3776, 8192,
  1, 28, 3776, 8192,
  1, 12, 3776, 8192,
  1, 12, 3776, 8192,
  1, 12, 3776, 8192,
  1, 0, 188, 8192,
  1, 12, 3776, 8192,
  1, 12, 3804, 8192,
  1, 12, 3804, 8192,
  1, 12, 3776, 8192,
  1, 0, 180, 8192,
  1, 12, 3792, 8192,
  1, 12, 3792, 8192,
  1, 12, 3792, 8192,
  1, 0, 156, 8192,
  1, 0, 156, 8192,
  1, 0, 176, 8192,
  0, 0, 160, 8192,
  0, 0, 160, 8192,
  0, 0, 128, 8192,
  0, 0, 128, 8192,
  0, 0, 128, 8192,
  0, 0, 128, 8192,
  0, 0, 128, 8192,
  0, 0, 128, 8192,
  0, 0, 128, 8192,
  0, 0, 128, 8192,
  0, 0, 128, 8192,
  0, 0, 160, 8192,
  0, 0, 160, 8192,
  1, 0, 176, 8192,
  1, 0, 16, 4096,
  0, 0, 128, 0,
  0, 0, 128, 0,
  0, 0, 128, 0,
  0, 0, 160, 8192,
  0, 0, 160, 8192,
  0, 0, 160, 8192,
  0, 0, 160, 8192,
  0, 0, 160, 8192,
  0, 0, 160, 8192,
  0, 0, 160, 8192,
  0, 0, 160, 8192,
  0, 0, 128, 0,
  1, 0, 144, 0,
  0, 0, 128, 0,
  0, 0, 128, 0,
  0, 0, 128, 0,
  0, 0, 128, 0,
  0, 0, 0, 4096,
  0, 0, 0, 4096,
  0, 0, 0, 4096,
  1, 0, 16, 4096,
  1, 0, 144, 8192,
  1, 0, 144, 8192,
  1, 0, 144, 8192,
  0, 0, 128, 8192,
  1, 0, 144, 8192,
  1, 0, 144, 8192,
  1, 0, 144, 8192,
  1, 0, 144, 8192,
  0, 0, 128, 8192,
  1, 0, 144, 8192,
  0, 0, 128, 8192,
  1, 0, 144, 8192,
  1, 0, 144, 8192,
  0, 0, 128, 8192,
  0, 0, 128, 8192,
  0, 0, 128, 8192,
  0, 0, 128, 8192,
  0, 0, 128, 8192,
  0, 0, 128, 8192,
  0, 0, 128, 8192,
  1, 0, 172, 8192,
  0, 0, 160, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  0, 0, 160, 8192,
  1, 0, 172, 8192,
  1, 0, 188, 8192,
  1, 0, 180, 8192,
  1, 0, 188, 8192,
  1, 0, 180, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  0, 0, 160, 8192,
  0, 0, 160, 8192,
  0, 0, 160, 8192,
  0, 0, 160, 8192,
  0, 0, 160, 8192,
  1, 12, 3776, 8192,
  0, 0, 160, 8192,
  0, 0, 160, 8192,
  1, 12, 3776, 8192,
  1, 0, 176, 8192,
  0, 0, 160, 8192,
  1, 0, 180, 8192,
  1, 12, 3804, 8192,
  1, 12, 3776, 8192,
  1, 12, 3792, 8192,
  1, 12, 3792, 8192,
  1, 12, 3792, 8192,
  1, 12, 3792, 8192,
  1, 0, 156, 8192,
  1, 0, 156, 8192,
  1, 0, 180, 8192,
  0, 0, 160, 8192,
  0, 0, 160, 8192,
  0, 0, 128, 8192,
  0, 0, 128, 8192,
  0, 0, 128, 8192,
  0, 0, 128, 8192,
  0, 0, 128, 8192,
  0, 0, 128, 8192,
  0, 0, 160, 8192,
  0, 0, 160, 8192,
  0, 0, 160, 8192,
  1, 0, 176, 8192,
  1, 0, 176, 8192,
  1, 0, 176, 8192,
  1, 0, 16, 4096,
  0, 0, 128, 0,
  0, 0, 128, 0,
  1, 0, 144, 8192,
  0, 0, 160, 8192,
  0, 0, 160, 8192,
  0, 0, 160, 8192,
  1, 0, 176, 8192,
  1, 0, 176, 8192,
  0, 0, 160, 8192,
  0, 0, 160, 8192,
  0, 0, 0, 4096,
  0, 0, 128, 0,
  0, 0, 128, 0,
  0, 0, 128, 0,
  0, 0, 128, 0,
  0, 0, 128, 0,
  0, 0, 128, 0,
  0, 0, 0, 4096,
  0, 0, 0, 4096,
  0, 0, 0, 4096,
  0, 0, 0, 4096,
  1, 0, 144, 8192,
  1, 0, 144, 8192,
  1, 0, 144, 8192,
  1, 0, 144, 8192,
  1, 0, 144, 8192,
  1, 0, 144, 8192,
  1, 0, 144, 8192,
  1, 0, 144, 8192,
  1, 0, 144, 8192,
  1, 0, 144, 8192,
  1, 0, 144, 8192,
  1, 0, 144, 8192,
  1, 0, 144, 8192,
  0, 0, 128, 8192,
  0, 0, 128, 8192,
  0, 0, 128, 8192,
  1, 0, 172, 8192,
  1, 0, 172, 8192,
  1, 0, 172, 8192,
  1, 0, 172, 8192,
  1, 0, 172, 8192,
  1, 0, 172, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  0, 0, 160, 8192,
  0, 0, 160, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 180, 8192,
  1, 0, 180, 8192,
  1, 28, 3776, 8192,
  1, 0, 176, 8192,
  0, 0, 160, 8192,
  1, 12, 3776, 8192,
  1, 12, 3776, 8192,
  1, 0, 180, 8192,
  0, 0, 160, 8192,
  1, 0, 188, 8192,
  1, 12, 3776, 8192,
  1, 12, 3776, 8192,
  1, 0, 188, 8192,
  1, 0, 180, 8192,
  1, 0, 188, 8192,
  1, 12, 3776, 8192,
  1, 12, 3792, 8192,
  1, 12, 3792, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 148, 8192,
  1, 0, 176, 8192,
  0, 0, 160, 8192,
  0, 0, 128, 8192,
  0, 0, 128, 8192,
  0, 0, 128, 8192,
  0, 0, 128, 8192,
  0, 0, 160, 8192,
  0, 0, 160, 8192,
  0, 0, 160, 8192,
  0, 0, 160, 8192,
  1, 0, 176, 8192,
  1, 0, 176, 8192,
  1, 0, 176, 8192,
  1, 0, 176, 8192,
  1, 0, 176, 8192,
  1, 0, 144, 8192,
  0, 0, 128, 0,
  0, 0, 128, 0,
  0, 0, 160, 8192,
  0, 0, 160, 8192,
  0, 0, 160, 8192,
  1, 0, 16, 4096,
  0, 0, 0, 4096,
  0, 0, 0, 4096,
  0, 0, 128, 0,
  0, 0, 128, 0,
  0, 0, 128, 0,
  1, 0, 144, 0,
  0, 0, 128, 0,
  0, 0, 128, 0,
  0, 0, 128, 0,
  0, 0, 128, 0,
  0, 0, 128, 0,
  0, 0, 128, 0,
  0, 0, 0, 4096,
  0, 0, 128, 0,
  1, 0, 144, 8192,
  1, 0, 144, 8192,
  1, 0, 144, 8192,
  1, 0, 144, 8192,
  0, 0, 128, 8192,
  1, 0, 144, 8192,
  1, 0, 144, 8192,
  1, 0, 144, 8192,
  1, 0, 144, 8192,
  1, 0, 144, 8192,
  1, 0, 148, 8192,
  1, 0, 144, 8192,
  0, 0, 128, 8192,
  0, 0, 128, 8192,
  0, 0, 128, 8192,
  1, 0, 172, 8192,
  1, 0, 172, 8192,
  0, 0, 160, 8192,
  0, 0, 160, 8192,
  1, 0, 172, 8192,
  1, 0, 172, 8192,
  1, 0, 172, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 172, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  0, 0, 160, 8192,
  1, 12, 3792, 8192,
  1, 12, 3776, 8192,
  1, 28, 3776, 8192,
  1, 28, 3776, 8192,
  1, 28, 3776, 8192,
  1, 12, 3776, 8192,
  1, 28, 3776, 8192,
  1, 12, 3776, 8192,
  1, 12, 3776, 8192,
  0, 0, 160, 8192,
  1, 12, 3776, 8192,
  1, 12, 3776, 8192,
  1, 0, 188, 8192,
  0, 0, 160, 8192,
  1, 12, 3776, 8192,
  1, 12, 3776, 8192,
  0, 0, 160, 8192,
  1, 12, 3776, 8192,
  1, 12, 3776, 8192,
  1, 12, 3776, 8192,
  0, 0, 160, 8192,
  1, 12, 3792, 8192,
  1, 12, 3792, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 176, 8192,
  1, 0, 176, 8192,
  0, 0, 160, 8192,
  0, 0, 128, 8192,
  0, 0, 128, 8192,
  0, 0, 160, 8192,
  0, 0, 160, 8192,
  0, 0, 160, 8192,
  0, 0, 160, 8192,
  0, 0, 160, 8192,
  1, 0, 176, 8192,
  1, 0, 176, 8192,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 176, 8192,
  1, 0, 176, 8192,
  1, 0, 176, 8192,
  1, 0, 180, 8192,
  1, 0, 16, 4096,
  0, 0, 160, 8192,
  0, 0, 160, 8192,
  0, 0, 160, 8192,
  1, 0, 16, 4096,
  0, 0, 128, 0,
  0, 0, 128, 0,
  0, 0, 128, 0,
  0, 0, 128, 0,
  0, 0, 128, 0,
  0, 0, 128, 0,
  0, 0, 128, 0,
  0, 0, 128, 0,
  0, 0, 128, 0,
  0, 0, 128, 0,
  0, 0, 128, 0,
  0, 0, 128, 0,
  0, 0, 128, 0,
  0, 0, 128, 0,
  1, 0, 144, 8192,
  1, 0, 144, 8192,
  1, 0, 144, 8192,
  0, 0, 128, 8192,
  1, 0, 144, 8192,
  1, 0, 144, 8192,
  1, 0, 144, 8192,
  0, 0, 128, 8192,
  1, 0, 144, 8192,
  1, 0, 144, 8192,
  1, 0, 144, 8192,
  0, 0, 128, 8192,
  0, 0, 128, 8192,
  0, 0, 128, 8192,
  0, 0, 128, 8192,
  1, 0, 172, 8192,
  1, 0, 188, 8192,
  1, 0, 180, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 172, 8192,
  1, 0, 172, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 172, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 176, 8192,
  1, 12, 3792, 8192,
  1, 12, 3792, 8192,
  1, 12, 3792, 8192,
  1, 12, 3792, 8192,
  1, 12, 3776, 8192,
  1, 28, 3776, 8192,
  1, 0, 188, 8192,
  0, 0, 160, 8192,
  0, 0, 160, 8192,
  1, 12, 3776, 8192,
  1, 12, 3776, 8192,
  1, 12, 3776, 8192,
  1, 12, 3776, 8192,
  1, 12, 3776, 8192,
  1, 12, 3776, 8192,
  1, 12, 3776, 8192,
  1, 12, 3776, 8192,
  0, 0, 160, 8192,
  0, 0, 160, 8192,
  1, 0, 180, 8192,
  1, 0, 176, 8192,
  1, 0, 176, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 156, 8192,
  1, 0, 188, 8192,
  1, 0, 176, 8192,
  1, 0, 144, 8192,
  1, 0, 176, 8192,
  0, 0, 160, 8192,
  0, 0, 160, 8192,
  0, 0, 160, 8192,
  0, 0, 160, 8192,
  0, 0, 160, 8192,
  0, 0, 160, 8192,
  0, 0, 160, 8192,
  1, 0, 176, 8192,
  1, 0, 176, 8192,
  1, 0, 16, 4096,
  0, 0, 128, 0,
  0, 0, 128, 0,
  1, 0, 16, 4096,
  1, 0, 176, 8192,
  1, 0, 176, 8192,
  1, 0, 48, 4096,
  1, 0, 16, 4096,
  1, 0, 144, 8192,
  1, 0, 48, 4096,
  1, 0, 16, 4096,
  0, 0, 128, 0,
  0, 0, 128, 0,
  0, 0, 128, 0,
  0, 0, 128, 0,
  0, 0, 128, 0,
  0, 0, 128, 0,
  0, 0, 128, 0,
  0, 0, 128, 0,
  0, 0, 128, 0,
  0, 0, 128, 0,
  0, 0, 128, 0,
  0, 0, 128, 0,
  0, 0, 128, 0,
  0, 0, 128, 0,
  0, 0, 128, 0,
  1, 0, 144, 8192,
  1, 0, 144, 8192,
  1, 0, 144, 8192,
  1, 0, 144, 8192,
  0, 0, 128, 8192,
  1, 0, 144, 8192,
  1, 0, 148, 8192,
  1, 0, 144, 8192,
  1, 0, 144, 8192,
  0, 0, 128, 8192,
  0, 0, 128, 8192,
  0, 0, 128, 8192,
  0, 0, 128, 8192,
  0, 0, 160, 8192,
  1, 0, 172, 8192,
  1, 0, 172, 8192,
  1, 0, 188, 8192,
  1, 0, 180, 8192,
  1, 0, 172, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 172, 8192,
  1, 0, 172, 8192,
  1, 0, 172, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 176, 8192,
  1, 0, 176, 8192,
  1, 0, 188, 8192,
  1, 12, 3792, 8192,
  1, 12, 3792, 8192,
  1, 0, 180, 8192,
  1, 0, 180, 8192,
  1, 0, 172, 8192,
  0, 0, 160, 8192,
  1, 12, 3776, 8192,
  1, 12, 3776, 8192,
  1, 12, 3776, 8192,
  1, 12, 3776, 8192,
  1, 12, 3776, 8192,
  1, 12, 3776, 8192,
  1, 12, 3776, 8192,
  1, 12, 3776, 8192,
  1, 12, 3776, 8192,
  0, 0, 160, 8192,
  1, 0, 176, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 148, 8192,
  1, 0, 180, 8192,
  1, 0, 176, 8192,
  1, 0, 176, 8192,
  1, 0, 176, 8192,
  1, 0, 176, 8192,
  0, 0, 160, 8192,
  0, 0, 160, 8192,
  0, 0, 160, 8192,
  0, 0, 160, 8192,
  1, 0, 176, 8192,
  1, 0, 176, 8192,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 144, 0,
  0, 0, 128, 0,
  0, 0, 128, 0,
  1, 0, 16, 4096,
  1, 0, 48, 4096,
  1, 0, 48, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  0, 0, 0, 4096,
  0, 0, 128, 0,
  1, 0, 16, 4096,
  0, 0, 0, 4096,
  0, 0, 128, 0,
  0, 0, 128, 0,
  0, 0, 128, 0,
  0, 0, 128, 0,
  0, 0, 128, 0,
  0, 0, 128, 0,
  0, 0, 128, 0,
  0, 0, 128, 0,
  0, 0, 128, 0,
  0, 0, 128, 0,
  1, 0, 144, 8192,
  1, 0, 144, 8192,
  1, 0, 144, 8192,
  1, 0, 144, 8192,
  1, 0, 144, 8192,
  1, 0, 144, 8192,
  1, 0, 144, 8192,
  1, 0, 144, 8192,
  1, 0, 144, 8192,
  1, 0, 144, 8192,
  0, 0, 128, 8192,
  0, 0, 128, 8192,
  0, 0, 128, 8192,
  1, 0, 172, 8192,
  1, 0, 172, 8192,
  1, 0, 188, 8192,
  0, 0, 160, 8192,
  0, 0, 160, 8192,
  1, 0, 172, 8192,
  1, 0, 172, 8192,
  1, 0, 172, 8192,
  1, 0, 188, 8192,
  1, 0, 140, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 164, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 180, 8192,
  1, 0, 180, 8192,
  1, 0, 176, 8192,
  1, 0, 176, 8192,
  1, 0, 180, 8192,
  1, 0, 188, 8192,
  1, 0, 164, 8192,
  1, 0, 188, 8192,
  0, 0, 160, 8192,
  1, 12, 3776, 8192,
  1, 12, 3776, 8192,
  1, 12, 3776, 8192,
  1, 12, 3776, 8192,
  1, 12, 3776, 8192,
  1, 12, 3776, 8192,
  1, 12, 3776, 8192,
  1, 12, 3776, 8192,
  1, 0, 180, 8192,
  1, 0, 188, 8192,
  1, 12, 3792, 8192,
  1, 0, 156, 8192,
  1, 0, 156, 8192,
  1, 0, 176, 8192,
  1, 0, 176, 8192,
  1, 0, 176, 8192,
  1, 0, 176, 8192,
  1, 0, 180, 8192,
  1, 0, 176, 8192,
  1, 0, 48, 4096,
  1, 0, 176, 8192,
  1, 0, 176, 8192,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  0, 0, 0, 4096,
  0, 0, 0, 4096,
  0, 0, 0, 4096,
  0, 0, 128, 0,
  0, 0, 128, 0,
  0, 0, 128, 0,
  1, 0, 144, 0,
  0, 0, 128, 0,
  0, 0, 128, 0,
  0, 0, 128, 0,
  0, 0, 128, 0,
  0, 0, 128, 0,
  0, 0, 128, 0,
  0, 0, 128, 0,
  1, 0, 144, 8192,
  1, 0, 144, 8192,
  1, 0, 144, 8192,
  1, 0, 144, 8192,
  1, 0, 144, 8192,
  1, 0, 144, 8192,
  1, 0, 144, 8192,
  1, 0, 144, 8192,
  0, 0, 128, 8192,
  0, 0, 128, 8192,
  0, 0, 128, 8192,
  0, 0, 128, 8192,
  1, 0, 172, 8192,
  1, 0, 172, 8192,
  0, 0, 160, 8192,
  1, 12, 3776, 8192,
  1, 12, 3776, 8192,
  0, 0, 160, 8192,
  0, 0, 160, 8192,
  1, 0, 172, 8192,
  1, 0, 172, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 12, 3792, 8192,
  1, 12, 3792, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  0, 0, 160, 8192,
  0, 0, 160, 8192,
  1, 12, 3776, 8192,
  1, 12, 3776, 8192,
  1, 0, 188, 8192,
  1, 12, 3776, 8192,
  1, 12, 3776, 8192,
  1, 12, 3776, 8192,
  1, 0, 176, 8192,
  1, 0, 188, 8192,
  1, 12, 3792, 8192,
  1, 0, 156, 8192,
  1, 0, 156, 8192,
  1, 0, 156, 8192,
  1, 0, 176, 8192,
  1, 0, 176, 8192,
  1, 0, 176, 8192,
  1, 0, 176, 8192,
  1, 0, 188, 8192,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 144, 0,
  0, 0, 128, 0,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 48, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  0, 0, 128, 0,
  0, 0, 128, 0,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  0, 0, 0, 4096,
  0, 0, 0, 4096,
  0, 0, 0, 4096,
  0, 0, 128, 0,
  0, 0, 128, 0,
  0, 0, 128, 8192,
  0, 0, 128, 8192,
  0, 0, 128, 8192,
  0, 0, 128, 0,
  0, 0, 32, 4096,
  0, 0, 128, 0,
  0, 0, 128, 0,
  0, 0, 128, 0,
  0, 0, 128, 0,
  1, 0, 144, 8192,
  1, 0, 144, 8192,
  1, 0, 144, 8192,
  1, 0, 144, 8192,
  1, 0, 144, 8192,
  1, 0, 144, 8192,
  1, 0, 144, 8192,
  0, 0, 128, 8192,
  0, 0, 128, 8192,
  0, 0, 128, 8192,
  0, 0, 128, 8192,
  1, 0, 172, 8192,
  1, 0, 172, 8192,
  1, 0, 188, 8192,
  0, 0, 160, 8192,
  1, 12, 3776, 8192,
  1, 12, 3780, 8192,
  1, 0, 164, 8192,
  1, 0, 172, 8192,
  1, 0, 172, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  0, 0, 160, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 12, 3792, 8192,
  1, 0, 188, 8192,
  1, 0, 176, 8192,
  1, 0, 176, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 12, 3776, 8192,
  1, 12, 3776, 8192,
  1, 12, 3776, 8192,
  1, 12, 3776, 8192,
  1, 0, 176, 8192,
  0, 0, 160, 8192,
  1, 12, 3792, 8192,
  1, 12, 3792, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 176, 8192,
  1, 0, 176, 8192,
  1, 0, 176, 8192,
  1, 0, 188, 8192,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 48, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 48, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  0, 0, 32, 4096,
  1, 0, 144, 0,
  0, 0, 128, 0,
  1, 0, 144, 0,
  0, 0, 128, 0,
  0, 0, 128, 8192,
  0, 0, 160, 8192,
  0, 0, 160, 8192,
  0, 0, 32, 4096,
  0, 0, 32, 4096,
  0, 0, 128, 0,
  0, 0, 128, 0,
  0, 0, 128, 0,
  1, 0, 144, 8192,
  1, 0, 144, 8192,
  1, 0, 148, 8192,
  1, 0, 144, 8192,
  1, 0, 148, 8192,
  1, 0, 144, 8192,
  0, 0, 128, 8192,
  0, 0, 128, 8192,
  0, 0, 128, 8192,
  0, 0, 128, 8192,
  1, 0, 172, 8192,
  1, 12, 3776, 8192,
  1, 12, 3788, 8192,
  1, 12, 3788, 8192,
  1, 12, 3776, 8192,
  1, 0, 180, 8192,
  1, 12, 3776, 8192,
  1, 0, 172, 8192,
  1, 0, 172, 8192,
  0, 0, 160, 8192,
  1, 0, 164, 8192,
  1, 0, 164, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 180, 8192,
  1, 0, 180, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 12, 3792, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 156, 8192,
  1, 12, 3776, 8192,
  1, 12, 3776, 8192,
  1, 12, 3776, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 188, 8192,
  1, 0, 176, 8192,
  1, 0, 176, 8192,
  1, 0, 180, 8192,
  1, 0, 188, 8192,
  1, 0, 144, 0,
  1, 0, 144, 0,
  1, 0, 16, 4096,
  1, 0, 48, 4096,
  1, 0, 48, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 48, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 16, 4096,
  1, 0, 48, 4096,
  1, 0, 16, 4096,
  1, 0, 48, 4096,
  1, 0, 48, 4096,
  0, 0, 32, 4096,
  1, 0, 144, 0,
  1, 0, 144, 0,
  1, 0, 144, 0,
  0, 0, 32, 4096,
  0, 0, 160, 8192,
  0, 0, 160, 8192,
  0, 0, 128, 0,
  0, 0, 32, 4096,
  0, 0, 128, 0,
  1, 0, 144, 0,
  1, 0, 16, 4096 ;

 RAzi_angle =
  46.83, 47.63, 48.37, 49.08, 49.75, 50.39, 50.99, 51.57, 52.12, 52.66, 
    53.18, 53.67, 54.14, 54.61, 55.07, 55.51, 55.94, 56.35, 56.76, 57.16, 
    57.55, 57.93, 58.3, 58.67, 59.03, 59.39, 59.73, 60.07, 60.41, 60.75, 
    61.08, 61.4, 61.72, 62.04, 62.36, 62.68, 62.99, 63.29, 63.59, 63.89, 
    64.18, 64.46, 64.73, 64.98, 65.19, 65.31, 65.16, 63.13, -110.08, -111.78, 
    -111.87, -111.73, -111.5, -111.23, -110.93, -110.62, -110.31, -109.98, 
    -109.64, -109.29, -108.94, -108.58, -108.21, -107.82, -107.43, -107.04, 
    -106.64, -106.22, -105.79, -105.35, -104.9, -104.44, -103.97, -103.48, 
    -102.96, -102.44, -101.9, -101.34, -100.75, -100.14, -99.51, -98.85, 
    -98.16, -97.42, -96.65, -95.85, -95.02, -94.13, -93.17, -92.14, -91.06, 
    -89.91, -88.67, -87.31, -85.83, -84.24,
  46.59, 47.39, 48.15, 48.86, 49.53, 50.15, 50.76, 51.34, 51.91, 52.44, 
    52.95, 53.45, 53.94, 54.41, 54.86, 55.3, 55.73, 56.15, 56.56, 56.96, 
    57.34, 57.72, 58.11, 58.48, 58.84, 59.19, 59.54, 59.89, 60.23, 60.57, 
    60.89, 61.22, 61.55, 61.87, 62.19, 62.5, 62.81, 63.12, 63.43, 63.72, 
    64.01, 64.29, 64.57, 64.82, 65.02, 65.14, 65, 62.83, -110.27, -111.92, 
    -112.01, -111.87, -111.63, -111.36, -111.07, -110.76, -110.44, -110.1, 
    -109.76, -109.42, -109.06, -108.7, -108.32, -107.93, -107.55, -107.15, 
    -106.74, -106.32, -105.89, -105.45, -105, -104.54, -104.05, -103.56, 
    -103.05, -102.53, -101.97, -101.4, -100.81, -100.2, -99.57, -98.9, 
    -98.19, -97.45, -96.69, -95.89, -95.03, -94.12, -93.16, -92.15, -91.06, 
    -89.88, -88.61, -87.26, -85.79, -84.19,
  46.36, 47.18, 47.93, 48.63, 49.3, 49.94, 50.55, 51.13, 51.69, 52.22, 52.74, 
    53.25, 53.73, 54.2, 54.65, 55.09, 55.53, 55.95, 56.35, 56.75, 57.14, 
    57.53, 57.91, 58.28, 58.64, 59, 59.35, 59.7, 60.04, 60.38, 60.71, 61.05, 
    61.37, 61.69, 62.01, 62.33, 62.64, 62.95, 63.25, 63.55, 63.85, 64.13, 
    64.41, 64.65, 64.87, 64.99, 64.85, 62.76, -110.38, -112.08, -112.17, 
    -112.02, -111.78, -111.51, -111.22, -110.9, -110.57, -110.24, -109.9, 
    -109.55, -109.19, -108.82, -108.44, -108.06, -107.67, -107.26, -106.85, 
    -106.43, -106, -105.56, -105.09, -104.62, -104.15, -103.65, -103.14, 
    -102.6, -102.04, -101.47, -100.88, -100.26, -99.61, -98.93, -98.23, 
    -97.5, -96.72, -95.9, -95.04, -94.14, -93.18, -92.14, -91.02, -89.84, 
    -88.59, -87.23, -85.73, -84.08,
  46.15, 46.95, 47.7, 48.41, 49.08, 49.72, 50.33, 50.91, 51.47, 52.02, 52.53, 
    53.03, 53.51, 53.98, 54.44, 54.89, 55.32, 55.74, 56.15, 56.55, 56.95, 
    57.33, 57.7, 58.08, 58.45, 58.81, 59.16, 59.5, 59.85, 60.19, 60.53, 
    60.86, 61.18, 61.51, 61.83, 62.15, 62.46, 62.77, 63.08, 63.38, 63.68, 
    63.96, 64.23, 64.49, 64.7, 64.83, 64.69, 62.64, -110.54, -112.23, 
    -112.32, -112.16, -111.93, -111.65, -111.35, -111.04, -110.71, -110.38, 
    -110.03, -109.67, -109.31, -108.95, -108.57, -108.18, -107.78, -107.37, 
    -106.97, -106.54, -106.1, -105.65, -105.19, -104.72, -104.24, -103.73, 
    -103.21, -102.67, -102.12, -101.54, -100.94, -100.31, -99.67, -99, 
    -98.29, -97.53, -96.74, -95.92, -95.07, -94.15, -93.17, -92.12, -91.02, 
    -89.84, -88.56, -87.16, -85.65, -84.01,
  45.91, 46.71, 47.48, 48.19, 48.86, 49.49, 50.1, 50.69, 51.25, 51.79, 52.31, 
    52.81, 53.3, 53.77, 54.23, 54.67, 55.11, 55.53, 55.95, 56.35, 56.74, 
    57.12, 57.51, 57.89, 58.25, 58.61, 58.96, 59.31, 59.66, 60, 60.34, 60.67, 
    61, 61.32, 61.64, 61.96, 62.28, 62.6, 62.91, 63.21, 63.5, 63.79, 64.07, 
    64.32, 64.53, 64.66, 64.52, 62.33, -110.72, -112.37, -112.46, -112.31, 
    -112.07, -111.79, -111.49, -111.18, -110.85, -110.51, -110.16, -109.81, 
    -109.45, -109.07, -108.68, -108.29, -107.9, -107.5, -107.07, -106.64, 
    -106.2, -105.75, -105.29, -104.81, -104.32, -103.82, -103.3, -102.76, 
    -102.19, -101.6, -101, -100.38, -99.73, -99.04, -98.31, -97.56, -96.78, 
    -95.96, -95.08, -94.15, -93.16, -92.12, -91, -89.79, -88.49, -87.11, 
    -85.61, -83.96,
  45.68, 46.5, 47.25, 47.95, 48.62, 49.26, 49.88, 50.47, 51.02, 51.56, 52.09, 
    52.6, 53.08, 53.55, 54.01, 54.46, 54.9, 55.32, 55.73, 56.13, 56.53, 
    56.93, 57.31, 57.68, 58.04, 58.41, 58.77, 59.12, 59.46, 59.81, 60.15, 
    60.48, 60.81, 61.13, 61.46, 61.78, 62.11, 62.42, 62.72, 63.03, 63.33, 
    63.62, 63.9, 64.15, 64.37, 64.5, 64.35, 62.24, -110.82, -112.53, -112.62, 
    -112.46, -112.22, -111.95, -111.65, -111.32, -110.99, -110.65, -110.3, 
    -109.94, -109.57, -109.2, -108.82, -108.43, -108.02, -107.61, -107.19, 
    -106.76, -106.32, -105.86, -105.39, -104.91, -104.42, -103.91, -103.38, 
    -102.83, -102.26, -101.69, -101.08, -100.44, -99.77, -99.08, -98.37, 
    -97.62, -96.81, -95.97, -95.09, -94.17, -93.18, -92.12, -90.97, -89.76, 
    -88.48, -87.08, -85.54, -83.85,
  45.46, 46.26, 47.01, 47.72, 48.4, 49.04, 49.65, 50.23, 50.8, 51.35, 51.87, 
    52.37, 52.86, 53.33, 53.8, 54.25, 54.68, 55.1, 55.52, 55.93, 56.33, 
    56.71, 57.1, 57.48, 57.85, 58.21, 58.57, 58.92, 59.27, 59.62, 59.95, 
    60.29, 60.62, 60.95, 61.28, 61.6, 61.92, 62.23, 62.55, 62.85, 63.15, 
    63.44, 63.72, 63.98, 64.2, 64.33, 64.19, 62.12, -111.02, -112.69, 
    -112.77, -112.62, -112.38, -112.09, -111.78, -111.47, -111.13, -110.79, 
    -110.43, -110.07, -109.71, -109.33, -108.94, -108.54, -108.14, -107.73, 
    -107.31, -106.87, -106.42, -105.96, -105.5, -105.02, -104.52, -104, 
    -103.46, -102.92, -102.35, -101.75, -101.13, -100.5, -99.84, -99.15, 
    -98.42, -97.65, -96.84, -96, -95.12, -94.17, -93.16, -92.09, -90.96, 
    -89.75, -88.44, -87.01, -85.46, -83.79,
  45.21, 46.02, 46.78, 47.49, 48.16, 48.8, 49.41, 50.01, 50.58, 51.12, 51.64, 
    52.15, 52.64, 53.12, 53.58, 54.02, 54.46, 54.9, 55.31, 55.72, 56.11, 
    56.51, 56.9, 57.27, 57.64, 58, 58.36, 58.72, 59.08, 59.42, 59.76, 60.1, 
    60.43, 60.76, 61.09, 61.41, 61.74, 62.06, 62.37, 62.67, 62.97, 63.27, 
    63.55, 63.82, 64.03, 64.17, 64.04, 61.88, -111.26, -112.87, -112.94, 
    -112.78, -112.53, -112.25, -111.95, -111.62, -111.28, -110.93, -110.58, 
    -110.22, -109.85, -109.46, -109.07, -108.67, -108.27, -107.85, -107.42, 
    -106.98, -106.54, -106.08, -105.6, -105.11, -104.6, -104.09, -103.56, 
    -103.01, -102.42, -101.82, -101.21, -100.57, -99.9, -99.19, -98.45, 
    -97.69, -96.89, -96.04, -95.12, -94.17, -93.17, -92.1, -90.95, -89.7, 
    -88.38, -86.96, -85.42, -83.72,
  44.97, 45.79, 46.54, 47.25, 47.92, 48.57, 49.19, 49.78, 50.34, 50.88, 
    51.42, 51.93, 52.42, 52.89, 53.35, 53.81, 54.25, 54.68, 55.09, 55.5, 
    55.91, 56.3, 56.68, 57.06, 57.43, 57.8, 58.17, 58.52, 58.87, 59.22, 
    59.56, 59.91, 60.24, 60.57, 60.9, 61.23, 61.55, 61.87, 62.18, 62.49, 
    62.8, 63.1, 63.38, 63.64, 63.87, 64, 63.88, 61.81, -111.34, -113.04, 
    -113.11, -112.94, -112.7, -112.41, -112.1, -111.77, -111.43, -111.08, 
    -110.73, -110.36, -109.98, -109.59, -109.21, -108.81, -108.39, -107.97, 
    -107.54, -107.11, -106.65, -106.18, -105.7, -105.21, -104.71, -104.19, 
    -103.65, -103.08, -102.5, -101.91, -101.28, -100.63, -99.95, -99.25, 
    -98.51, -97.74, -96.91, -96.04, -95.15, -94.2, -93.18, -92.09, -90.92, 
    -89.68, -88.36, -86.92, -85.33, -83.61,
  44.74, 45.55, 46.31, 47.03, 47.71, 48.35, 48.96, 49.55, 50.12, 50.67, 
    51.19, 51.69, 52.18, 52.67, 53.14, 53.59, 54.02, 54.45, 54.88, 55.29, 
    55.69, 56.08, 56.47, 56.85, 57.23, 57.6, 57.95, 58.31, 58.67, 59.02, 
    59.36, 59.7, 60.04, 60.37, 60.71, 61.03, 61.36, 61.68, 62, 62.31, 62.61, 
    62.91, 63.19, 63.46, 63.69, 63.83, 63.7, 61.65, -111.58, -113.2, -113.27, 
    -113.1, -112.85, -112.56, -112.25, -111.92, -111.58, -111.23, -110.86, 
    -110.5, -110.12, -109.74, -109.34, -108.93, -108.52, -108.1, -107.67, 
    -107.22, -106.76, -106.29, -105.82, -105.32, -104.81, -104.28, -103.74, 
    -103.18, -102.59, -101.98, -101.34, -100.69, -100.02, -99.31, -98.56, 
    -97.76, -96.94, -96.09, -95.18, -94.2, -93.17, -92.08, -90.92, -89.67, 
    -88.3, -86.84, -85.27, -83.56,
  44.49, 45.31, 46.07, 46.79, 47.46, 48.1, 48.72, 49.31, 49.88, 50.42, 50.95, 
    51.47, 51.96, 52.44, 52.9, 53.36, 53.8, 54.24, 54.66, 55.06, 55.46, 
    55.87, 56.26, 56.64, 57.01, 57.38, 57.75, 58.11, 58.46, 58.81, 59.16, 
    59.5, 59.84, 60.17, 60.5, 60.83, 61.17, 61.49, 61.81, 62.12, 62.42, 
    62.73, 63.02, 63.28, 63.51, 63.65, 63.52, 61.37, -111.76, -113.36, 
    -113.43, -113.26, -113.01, -112.73, -112.41, -112.08, -111.73, -111.37, 
    -111.01, -110.65, -110.27, -109.87, -109.47, -109.07, -108.65, -108.23, 
    -107.79, -107.34, -106.88, -106.41, -105.93, -105.42, -104.9, -104.38, 
    -103.84, -103.27, -102.67, -102.05, -101.42, -100.77, -100.08, -99.35, 
    -98.6, -97.82, -97, -96.11, -95.18, -94.21, -93.19, -92.08, -90.89, 
    -89.61, -88.26, -86.81, -85.22, -83.46,
  44.26, 45.08, 45.83, 46.54, 47.22, 47.87, 48.48, 49.07, 49.64, 50.19, 
    50.73, 51.24, 51.73, 52.2, 52.68, 53.14, 53.58, 54.01, 54.43, 54.84, 
    55.25, 55.65, 56.04, 56.42, 56.8, 57.17, 57.54, 57.9, 58.25, 58.61, 
    58.96, 59.3, 59.64, 59.97, 60.31, 60.65, 60.97, 61.29, 61.61, 61.93, 
    62.24, 62.54, 62.83, 63.1, 63.33, 63.48, 63.36, 61.36, -111.9, -113.55, 
    -113.61, -113.44, -113.19, -112.89, -112.57, -112.23, -111.89, -111.53, 
    -111.17, -110.79, -110.41, -110.02, -109.62, -109.21, -108.78, -108.35, 
    -107.92, -107.47, -107.01, -106.52, -106.03, -105.53, -105.02, -104.49, 
    -103.93, -103.35, -102.76, -102.15, -101.5, -100.83, -100.14, -99.42, 
    -98.67, -97.87, -97.02, -96.14, -95.21, -94.23, -93.18, -92.06, -90.86, 
    -89.6, -88.25, -86.75, -85.12, -83.36 ;

 RFlag =
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888 ;

 RR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 13, 20, 13, 11, 12, 9, 8, 0, 0, 
    6, 9, 0, 5, 7, 15, 16, 18, 13, 6, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, _, _, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 9, 13, 15, 32, 44, 31, 7, 16, 26, 23, 
    32, 34, 31, 24, 16, 14, 20, 16, 22, 24, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, 
    _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 6, 9, 12, 10, 9, 11, 9, 12, 12, 17, 13, 15, 16, 9, 14, 16, 
    13, 14, 14, 31, 16, 20, 20, 17, 34, 18, 14, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, 
    _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 5, 0, 6, 11, 10, 18, 12, 13, 11, 12, 8, 9, 12, 11, 11, 10, 6, 9, 13, 
    8, 11, 13, 8, 11, 18, 17, 17, 16, 14, 9, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, _, _, _, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, 
    _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 7, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 5, 12, 11, 9, 10, 19, 22, 19, 16, 16, 13, 12, 11, 12, 15, 15, 
    11, 15, 12, 12, 8, 13, 16, 12, 11, 9, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 18, 17, 9, 0, 0, 0, 0, 
    0, 0, 0, 6, 6, 6, 9, 11, 13, 15, 16, 16, 14, 15, 17, 15, 14, 11, 15, 11, 
    0, 15, 13, 16, 17, 12, 14, 12, 5, 7, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, _, _, 0, 0, 0, 0, _, 0, 0, 0, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 19, 13, 0, 0, 0, 0, 0, 
    0, 0, 5, 6, 0, 6, 10, 22, 15, 16, 16, 15, 15, 16, 33, 10, 8, 13, 14, 15, 
    15, 14, 15, 16, 14, 9, 14, 8, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, _, _, _, _, 0, 0, _, _, 0, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 0, 0, 0, 0, 0, 0, 0, 
    5, 10, 8, 6, 11, 13, 14, 21, 23, 19, 25, 16, 14, 16, 15, 17, 19, 16, 17, 
    15, 16, 15, 13, 10, 9, 11, 8, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 7, 0, 0, 0, 0, 0, 4, 0, 0, 
    0, 5, 6, 6, 9, 9, 8, 9, 9, 14, 11, 9, 13, 11, 9, 7, 12, 12, 14, 15, 13, 
    12, 11, 10, 10, 9, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, _, 0, 0, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 0, 0, _, _, _, 
    _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 7, 7, 7, 0, 0, 0, 0, 0, 0, 0, 
    0, 7, 0, 7, 6, 7, 5, 8, 9, 8, 10, 10, 10, 11, 8, 6, 5, 9, 16, 14, 12, 6, 
    10, 10, 10, 5, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 0, 0, 0, _, _, _, _, 
    _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 7, 9, 9, 8, 9, 0, 0, 0, 7, 12, 8, 
    6, 6, 5, 7, 6, 0, 7, 8, 9, 9, 12, 11, 11, 11, 16, 12, 7, 0, 0, 0, 0, 7, 
    7, 9, 10, 0, 5, 8, 7, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 0, 0, 0, _, _, _, 
    _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 8, 8, 6, 23, 7, 7, 0, 0, 0, 7, 10, 8, 
    6, 6, 0, 5, 5, 7, 13, 8, 8, 14, 10, 13, 9, 9, 8, 11, 8, 6, 0, 0, 0, 0, 0, 
    7, 9, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 0, 0, _, _, _, _, _ ;

 RWP =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, _, _, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 0, 0, 0, 0, 0, 
    0, 22, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, _, _, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 21, 0, 0, 17, 22, 18, 18, 
    19, 0, 16, 10, 13, 14, 0, 14, 11, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, _, _, _, _, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, 
    _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 0, 0, 16, 0, 
    0, 0, 14, 13, 13, 10, 7, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, _, _, _, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 0, 0, 16, 18, 0, 0, 0, 13, 
    13, 0, 0, 0, 11, 8, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, _, _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 16, 18, 20, 21, 20, 19, 23, 18, 18, 0, 15, 10, 0, 0, 
    12, 12, 0, 9, 14, 10, 0, 6, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, _, _, 0, 0, 0, 0, _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 15, 14, 17, 18, 17, 20, 0, 0, 0, 13, 14, 12, 11, 10, 
    9, 8, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    _, _, _, _, 0, 0, _, _, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 14, 0, 0, 0, 0, 12, 9, 10, 11, 10, 
    9, 8, 7, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 9, 8, 8, 7, 6, 
    6, 7, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, _, 0, 0, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 10, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 10, 0, 0, 0, 0, 0, 10, 9, 0, 7, 
    6, 8, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 0, 0, 0, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 10, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 0, 0, 0, 0, 0, 0, 0, 0, 5, 5, 6, 
    7, 0, 0, 7, 7, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 0, 0, 0, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 9, 9, 8, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 7, 
    6, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 0, 0, _, _, _, _, _ ;

 SFR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, _, _, _, _, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, _, _, _, _, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, _, _, _, _, _, _, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    _, _, _, _, _, _, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    _, _, _, _, _, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, 
    _, 0, _, _, _, _, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, 
    _, _, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, 0, 0, 0, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 0, _, _, _, _, _, _ ;

 SIce =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, 100, 100, _, _, _, _, _, _, _, _, _, _, 62, 58, 50, 38, 0, 0, 0, 0,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, 100, 100, _, _, _, _, _, _, _, _, _, 62, 58, 62, 52, 42, 0, 0, 
    0, 0,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, 0, 100, 100, 50, _, _, _, _, _, _, _, _, 62, 56, 58, 62, 56, 46, 0, 0, 
    0, 0,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, 0, 100, 100, _, _, _, _, _, _, _, _, 44, 52, 54, 58, 64, 62, 0, 38, 0, 
    0, 0,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, 38, 44, _, _, _, 0, 0, 40, 44, 44, 46, 58, 64, 64, 64, 0, 0, 0, 
    0, 0,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 100, 0, 
    _, _, _, _, 0, _, _, _, 36, 32, 32, 32, 38, 52, 60, 70, 76, 72, 0, 0, 0, 
    0, 0,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 100, 100, 
    100, 0, _, _, 0, 0, _, 0, 0, 22, 22, 24, 0, 42, 54, 62, 74, 78, 76, 0, 0, 
    0, 0, 0,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 0, 0, 100, 100, 
    100, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 46, 60, 66, 76, 80, 78, 70, 56, 
    0, 0, 0,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, 0, _, _, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 44, 56, 66, 72, _, _, 80, 72, 0, 48, 0, 0,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, 0, 0, 0, 98, 100, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 52, 64, 68, _, _, _, 80, 76, 66, 54, 
    46, 0,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 58, 68, 74, 78, _, _, _, 74, 72, 60, 0, 0,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, 100, 100, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 36, 54, 70, 76, 78, 76, _, _, 84, 76, 
    62, 0, 58 ;

 SIce_FY =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, 12, 96, _, _, _, _, _, _, _, _, _, _, 62, 58, 50, 38, 0, 0, 0, 0,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, 5, 76, _, _, _, _, _, _, _, _, _, 62, 58, 62, 52, 42, 0, 0, 0, 0,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, 0, 28, 18, 50, _, _, _, _, _, _, _, _, 62, 56, 58, 62, 56, 46, 0, 0, 
    0, 0,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, 0, 78, 86, _, _, _, _, _, _, _, _, 44, 52, 54, 58, 64, 62, 0, 38, 0, 
    0, 0,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, 38, 44, _, _, _, 0, 0, 37, 44, 44, 46, 58, 64, 64, 64, 0, 0, 0, 
    0, 0,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 100, 0, 
    _, _, _, _, 0, _, _, _, 31, 32, 32, 0, 38, 52, 60, 70, 76, 72, 0, 0, 0, 
    0, 0,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 100, 38, 
    86, 0, _, _, 0, 0, _, 0, 0, 0, 22, 24, 0, 42, 54, 62, 74, 78, 76, 0, 0, 
    0, 0, 0,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 0, 0, 100, 100, 
    100, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 46, 60, 66, 76, 80, 78, 70, 56, 
    0, 0, 0,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, 0, _, _, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 44, 56, 66, 72, _, _, 80, 72, 0, 48, 0, 0,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, 0, 0, 0, 98, 100, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 52, 64, 68, _, _, _, 80, 76, 66, 52, 
    45, 0,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 58, 68, 74, 78, _, _, _, 74, 72, 60, 0, 0,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, 100, 100, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 36, 54, 70, 76, 78, 76, _, _, 84, 76, 
    62, 0, 58 ;

 SIce_MY =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, 88, 4, _, _, _, _, _, _, _, _, _, _, 0, 0, 0, 0, 0, 0, 0, 0,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, 95, 24, _, _, _, _, _, _, _, _, _, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, 0, 72, 82, 0, _, _, _, _, _, _, _, _, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, 0, 22, 14, _, _, _, _, _, _, _, _, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, 0, 0, _, _, _, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 0, 0, 
    _, _, _, _, 0, _, _, _, 4, 0, 0, 31, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 0, 62, 14, 
    0, _, _, 0, 0, _, 0, 0, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, 0, _, _, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, 0, 0, 0, 0, 0, 0,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, 0, 0, 0, 1, 0, 0,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, 0, 0, 0, 0, 0,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, 0, 0, 0, 0, 0 ;

 SWE =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, _, _, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, _, _, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, _, _, _, _, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, _, _, _, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, _, _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, 
    0, 0, 0, 0, _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, 
    _, 0, 0, _, _, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, 0, 0, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 0, 0, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, 0, 0, 0, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 0, 0, 0, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 0, 0, _, _, _, _, _ ;

 SWP =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 SZ_angle =
  41.29, 41.39, 41.49, 41.59, 41.68, 41.78, 41.86, 41.95, 42.03, 42.11, 
    42.19, 42.27, 42.34, 42.41, 42.49, 42.56, 42.63, 42.69, 42.76, 42.82, 
    42.88, 42.95, 43.01, 43.07, 43.13, 43.18, 43.24, 43.3, 43.35, 43.41, 
    43.47, 43.52, 43.57, 43.63, 43.68, 43.74, 43.79, 43.84, 43.89, 43.95, 44, 
    44.05, 44.11, 44.16, 44.21, 44.27, 44.32, 44.37, 44.43, 44.48, 44.54, 
    44.59, 44.65, 44.7, 44.76, 44.82, 44.88, 44.94, 45, 45.06, 45.12, 45.18, 
    45.25, 45.31, 45.38, 45.45, 45.52, 45.59, 45.66, 45.74, 45.82, 45.9, 
    45.98, 46.06, 46.15, 46.24, 46.33, 46.43, 46.53, 46.64, 46.75, 46.86, 
    46.99, 47.11, 47.25, 47.39, 47.54, 47.7, 47.87, 48.06, 48.25, 48.47, 
    48.7, 48.95, 49.23, 49.54,
  41.44, 41.54, 41.64, 41.74, 41.83, 41.92, 42.01, 42.1, 42.18, 42.26, 42.34, 
    42.42, 42.49, 42.57, 42.64, 42.71, 42.77, 42.84, 42.91, 42.97, 43.03, 
    43.09, 43.16, 43.22, 43.28, 43.33, 43.39, 43.45, 43.5, 43.56, 43.61, 
    43.67, 43.72, 43.78, 43.83, 43.88, 43.94, 43.99, 44.04, 44.1, 44.15, 
    44.2, 44.25, 44.31, 44.36, 44.41, 44.46, 44.52, 44.57, 44.63, 44.68, 
    44.74, 44.79, 44.85, 44.91, 44.96, 45.02, 45.08, 45.14, 45.2, 45.26, 
    45.33, 45.39, 45.46, 45.52, 45.59, 45.66, 45.73, 45.81, 45.88, 45.96, 
    46.04, 46.12, 46.21, 46.29, 46.38, 46.48, 46.57, 46.68, 46.78, 46.89, 47, 
    47.13, 47.26, 47.39, 47.53, 47.68, 47.84, 48.01, 48.19, 48.39, 48.6, 
    48.83, 49.09, 49.36, 49.67,
  41.59, 41.69, 41.8, 41.89, 41.99, 42.08, 42.17, 42.25, 42.33, 42.41, 42.49, 
    42.57, 42.65, 42.72, 42.79, 42.86, 42.93, 42.99, 43.06, 43.12, 43.18, 
    43.25, 43.31, 43.37, 43.42, 43.48, 43.54, 43.6, 43.65, 43.71, 43.76, 
    43.82, 43.87, 43.92, 43.98, 44.03, 44.09, 44.14, 44.19, 44.24, 44.3, 
    44.35, 44.4, 44.45, 44.51, 44.56, 44.61, 44.67, 44.72, 44.77, 44.83, 
    44.88, 44.94, 45, 45.05, 45.11, 45.17, 45.23, 45.29, 45.35, 45.41, 45.47, 
    45.54, 45.6, 45.67, 45.74, 45.81, 45.88, 45.95, 46.02, 46.1, 46.18, 
    46.26, 46.35, 46.43, 46.52, 46.62, 46.71, 46.82, 46.92, 47.03, 47.15, 
    47.27, 47.39, 47.53, 47.67, 47.82, 47.98, 48.14, 48.33, 48.53, 48.74, 
    48.97, 49.22, 49.5, 49.81,
  41.74, 41.85, 41.95, 42.04, 42.14, 42.23, 42.32, 42.4, 42.49, 42.57, 42.65, 
    42.72, 42.79, 42.87, 42.94, 43.01, 43.08, 43.14, 43.21, 43.27, 43.33, 
    43.39, 43.45, 43.51, 43.57, 43.63, 43.69, 43.74, 43.8, 43.86, 43.91, 
    43.97, 44.02, 44.07, 44.13, 44.18, 44.23, 44.29, 44.34, 44.39, 44.44, 
    44.49, 44.55, 44.6, 44.65, 44.71, 44.76, 44.81, 44.87, 44.92, 44.98, 
    45.03, 45.08, 45.14, 45.2, 45.26, 45.31, 45.37, 45.43, 45.49, 45.55, 
    45.62, 45.68, 45.75, 45.81, 45.88, 45.95, 46.02, 46.09, 46.17, 46.25, 
    46.32, 46.4, 46.49, 46.58, 46.67, 46.76, 46.86, 46.96, 47.06, 47.17, 
    47.28, 47.4, 47.53, 47.67, 47.81, 47.95, 48.11, 48.28, 48.47, 48.66, 
    48.87, 49.1, 49.35, 49.63, 49.94,
  41.89, 42, 42.1, 42.2, 42.29, 42.38, 42.47, 42.55, 42.64, 42.72, 42.8, 
    42.87, 42.95, 43.02, 43.09, 43.16, 43.23, 43.29, 43.36, 43.42, 43.48, 
    43.54, 43.61, 43.67, 43.72, 43.78, 43.84, 43.89, 43.95, 44.01, 44.06, 
    44.11, 44.17, 44.22, 44.27, 44.33, 44.38, 44.43, 44.49, 44.54, 44.59, 
    44.64, 44.7, 44.75, 44.8, 44.85, 44.9, 44.96, 45.01, 45.07, 45.12, 45.18, 
    45.23, 45.29, 45.34, 45.4, 45.46, 45.52, 45.58, 45.64, 45.7, 45.76, 
    45.83, 45.89, 45.96, 46.02, 46.09, 46.16, 46.24, 46.31, 46.39, 46.47, 
    46.55, 46.63, 46.72, 46.81, 46.9, 47, 47.1, 47.2, 47.31, 47.43, 47.55, 
    47.67, 47.8, 47.94, 48.09, 48.25, 48.42, 48.6, 48.8, 49.01, 49.24, 49.49, 
    49.76, 50.07,
  42.04, 42.15, 42.25, 42.35, 42.44, 42.53, 42.62, 42.71, 42.79, 42.87, 
    42.95, 43.02, 43.1, 43.17, 43.24, 43.31, 43.38, 43.44, 43.51, 43.57, 
    43.63, 43.7, 43.76, 43.81, 43.87, 43.93, 43.99, 44.04, 44.1, 44.15, 
    44.21, 44.26, 44.32, 44.37, 44.42, 44.48, 44.53, 44.58, 44.63, 44.69, 
    44.74, 44.79, 44.84, 44.89, 44.95, 45, 45.05, 45.1, 45.16, 45.21, 45.27, 
    45.32, 45.38, 45.43, 45.49, 45.55, 45.6, 45.66, 45.72, 45.78, 45.84, 
    45.91, 45.97, 46.03, 46.1, 46.17, 46.24, 46.31, 46.38, 46.45, 46.53, 
    46.61, 46.69, 46.77, 46.86, 46.95, 47.04, 47.14, 47.24, 47.34, 47.45, 
    47.57, 47.69, 47.81, 47.94, 48.09, 48.23, 48.39, 48.56, 48.74, 48.93, 
    49.15, 49.37, 49.62, 49.9, 50.21,
  42.2, 42.3, 42.4, 42.5, 42.59, 42.68, 42.77, 42.86, 42.94, 43.02, 43.1, 
    43.17, 43.25, 43.32, 43.39, 43.46, 43.53, 43.59, 43.66, 43.72, 43.78, 
    43.84, 43.9, 43.96, 44.02, 44.08, 44.14, 44.19, 44.25, 44.3, 44.36, 
    44.41, 44.46, 44.52, 44.57, 44.62, 44.68, 44.73, 44.78, 44.83, 44.89, 
    44.94, 44.99, 45.04, 45.09, 45.15, 45.2, 45.25, 45.31, 45.36, 45.41, 
    45.47, 45.52, 45.58, 45.64, 45.69, 45.75, 45.81, 45.87, 45.93, 45.99, 
    46.05, 46.11, 46.18, 46.25, 46.31, 46.38, 46.45, 46.52, 46.6, 46.67, 
    46.75, 46.83, 46.92, 47, 47.09, 47.18, 47.28, 47.38, 47.48, 47.59, 47.7, 
    47.82, 47.95, 48.08, 48.22, 48.37, 48.53, 48.7, 48.88, 49.07, 49.28, 
    49.51, 49.76, 50.03, 50.33,
  42.35, 42.45, 42.55, 42.65, 42.74, 42.83, 42.92, 43.01, 43.09, 43.17, 
    43.25, 43.33, 43.4, 43.47, 43.54, 43.61, 43.68, 43.74, 43.81, 43.87, 
    43.93, 43.99, 44.06, 44.11, 44.17, 44.23, 44.29, 44.34, 44.4, 44.45, 
    44.51, 44.56, 44.61, 44.67, 44.72, 44.77, 44.83, 44.88, 44.93, 44.98, 
    45.03, 45.09, 45.14, 45.19, 45.24, 45.29, 45.35, 45.4, 45.45, 45.51, 
    45.56, 45.61, 45.67, 45.73, 45.78, 45.84, 45.9, 45.95, 46.01, 46.07, 
    46.13, 46.2, 46.26, 46.32, 46.39, 46.46, 46.52, 46.6, 46.67, 46.74, 
    46.82, 46.9, 46.98, 47.06, 47.14, 47.23, 47.33, 47.42, 47.52, 47.62, 
    47.73, 47.85, 47.97, 48.09, 48.22, 48.36, 48.51, 48.67, 48.83, 49.01, 
    49.21, 49.42, 49.64, 49.89, 50.16, 50.47,
  42.5, 42.61, 42.71, 42.8, 42.9, 42.99, 43.08, 43.16, 43.24, 43.32, 43.4, 
    43.48, 43.55, 43.62, 43.69, 43.76, 43.83, 43.89, 43.96, 44.02, 44.08, 
    44.15, 44.2, 44.26, 44.32, 44.38, 44.44, 44.49, 44.55, 44.6, 44.66, 
    44.71, 44.76, 44.82, 44.87, 44.92, 44.97, 45.03, 45.08, 45.13, 45.18, 
    45.23, 45.28, 45.34, 45.39, 45.44, 45.49, 45.55, 45.6, 45.65, 45.71, 
    45.76, 45.82, 45.87, 45.93, 45.98, 46.04, 46.1, 46.16, 46.22, 46.28, 
    46.34, 46.4, 46.47, 46.53, 46.6, 46.67, 46.74, 46.81, 46.88, 46.96, 
    47.04, 47.12, 47.2, 47.29, 47.38, 47.47, 47.56, 47.66, 47.77, 47.87, 
    47.99, 48.1, 48.23, 48.36, 48.5, 48.65, 48.8, 48.97, 49.15, 49.34, 49.55, 
    49.78, 50.02, 50.3, 50.61,
  42.65, 42.76, 42.86, 42.96, 43.05, 43.14, 43.23, 43.31, 43.4, 43.48, 43.55, 
    43.63, 43.7, 43.77, 43.84, 43.91, 43.98, 44.04, 44.11, 44.17, 44.23, 
    44.29, 44.35, 44.41, 44.47, 44.53, 44.58, 44.64, 44.7, 44.75, 44.8, 
    44.86, 44.91, 44.96, 45.02, 45.07, 45.12, 45.17, 45.23, 45.28, 45.33, 
    45.38, 45.43, 45.48, 45.54, 45.59, 45.64, 45.69, 45.75, 45.8, 45.85, 
    45.91, 45.96, 46.02, 46.07, 46.13, 46.19, 46.24, 46.3, 46.36, 46.42, 
    46.48, 46.55, 46.61, 46.68, 46.74, 46.81, 46.88, 46.95, 47.03, 47.1, 
    47.18, 47.26, 47.34, 47.43, 47.52, 47.61, 47.71, 47.81, 47.91, 48.01, 
    48.13, 48.25, 48.37, 48.5, 48.64, 48.78, 48.94, 49.11, 49.29, 49.48, 
    49.69, 49.91, 50.16, 50.43, 50.73,
  42.8, 42.91, 43.01, 43.11, 43.2, 43.29, 43.38, 43.46, 43.55, 43.63, 43.7, 
    43.78, 43.85, 43.93, 43.99, 44.06, 44.13, 44.2, 44.26, 44.32, 44.38, 
    44.44, 44.51, 44.56, 44.62, 44.68, 44.73, 44.79, 44.85, 44.9, 44.95, 
    45.01, 45.06, 45.11, 45.16, 45.22, 45.27, 45.32, 45.37, 45.42, 45.48, 
    45.53, 45.58, 45.63, 45.68, 45.73, 45.79, 45.84, 45.89, 45.95, 46, 46.05, 
    46.11, 46.16, 46.22, 46.27, 46.33, 46.39, 46.45, 46.51, 46.57, 46.63, 
    46.69, 46.76, 46.82, 46.89, 46.96, 47.03, 47.1, 47.17, 47.25, 47.33, 
    47.41, 47.49, 47.57, 47.66, 47.75, 47.85, 47.95, 48.05, 48.16, 48.27, 
    48.39, 48.51, 48.64, 48.78, 48.93, 49.08, 49.25, 49.42, 49.62, 49.83, 
    50.05, 50.29, 50.56, 50.87,
  42.96, 43.06, 43.16, 43.26, 43.35, 43.44, 43.53, 43.62, 43.7, 43.78, 43.86, 
    43.93, 44, 44.08, 44.15, 44.21, 44.28, 44.35, 44.41, 44.47, 44.53, 44.6, 
    44.65, 44.71, 44.77, 44.83, 44.88, 44.94, 44.99, 45.05, 45.1, 45.16, 
    45.21, 45.26, 45.31, 45.37, 45.42, 45.47, 45.52, 45.57, 45.62, 45.68, 
    45.73, 45.78, 45.83, 45.88, 45.93, 45.99, 46.04, 46.09, 46.15, 46.2, 
    46.25, 46.31, 46.37, 46.42, 46.48, 46.54, 46.59, 46.65, 46.71, 46.78, 
    46.84, 46.9, 46.97, 47.03, 47.1, 47.17, 47.24, 47.32, 47.39, 47.47, 
    47.55, 47.63, 47.71, 47.8, 47.89, 47.99, 48.09, 48.19, 48.3, 48.41, 
    48.52, 48.65, 48.78, 48.92, 49.06, 49.22, 49.38, 49.56, 49.76, 49.96, 
    50.18, 50.43, 50.7, 51.01 ;

 ScanTime_UTC = 5226.00048828125, 5229.00048828125, 5232.00048828125, 
    5234.00048828125, 5237.00048828125, 5240.00048828125, 5242.00048828125, 
    5245.00048828125, 5248.00048828125, 5250.00048828125, 5253.00048828125, 
    5256.00048828125 ;

 ScanTime_dom = 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30 ;

 ScanTime_doy = 181, 181, 181, 181, 181, 181, 181, 181, 181, 181, 181, 181 ;

 ScanTime_hour = 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1 ;

 ScanTime_minute = 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27 ;

 ScanTime_month = 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6 ;

 ScanTime_second = 6, 9, 12, 14, 17, 20, 22, 25, 28, 30, 33, 36 ;

 ScanTime_year = 2021, 2021, 2021, 2021, 2021, 2021, 2021, 2021, 2021, 2021, 
    2021, 2021 ;

 Sfc_type =
  2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 1, 1, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 1, 1, 1, 1, 0, 0, 0, 0,
  2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 1, 1, 2, 2, 2, 2, 2, 2, 2, 2, 2, 1, 1, 1, 1, 1, 0, 0, 0, 0,
  2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 0, 1, 1, 1, 2, 2, 2, 2, 2, 2, 2, 2, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0,
  2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 0, 1, 1, 2, 2, 2, 2, 2, 2, 2, 2, 1, 1, 1, 1, 1, 1, 0, 1, 0, 0, 0,
  2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 1, 1, 2, 2, 2, 0, 0, 1, 1, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0,
  2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 1, 0, 
    2, 2, 2, 2, 0, 2, 2, 2, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0,
  2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 1, 1, 1, 
    0, 2, 2, 0, 0, 2, 0, 0, 1, 1, 1, 0, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0,
  2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 0, 0, 1, 1, 1, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 1, 1, 0, 0, 0,
  2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 0, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 2, 2, 1, 1, 0, 1, 0, 0,
  2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 2, 2, 2, 1, 1, 1, 1, 1, 0,
  2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 2, 2, 2, 1, 1, 1, 0, 0,
  2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 2, 2, 1, 1, 1, 0, 1 ;

 Snow =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, _, _, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, _, _, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, _, _, _, _, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, _, _, _, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, _, _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, 
    0, 0, 0, 0, _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, 
    _, 0, 0, _, _, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, 0, 0, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 0, 0, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, 0, 0, 0, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 0, 0, 0, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 0, 0, _, _, _, _, _ ;

 SnowGS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, _, _, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, _, _, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, _, _, _, _, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, _, _, _, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, _, _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, 
    0, 0, 0, 0, _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, 
    _, 0, 0, _, _, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, 0, 0, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 0, 0, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, 0, 0, 0, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 0, 0, 0, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 0, 0, _, _, _, _, _ ;

 SurfM =
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888 ;

 SurfP =
  9620, 9332, 8760, 9070, 8653, 8316, 8488, 8747, 8906, 8985, 8700, 8896, 
    8499, 8956, 8856, 8638, 8345, 8958, 9325, 8754, 8589, 8933, 8842, 9413, 
    9838, 9781, 10002, 10018, 10018, 10018, 10010, 9885, 9936, 9831, 9905, 
    9862, 9855, 9930, 9781, 9912, 9971, 9853, 9890, 9870, 9858, 9909, 9801, 
    9755, 9796, 9822, 10007, 9900, 9652, 9721, 9939, 9974, 10018, 10027, 
    10027, 10018, 9968, 9912, 9708, 9924, 9862, 9756, 9560, 9441, 9480, 9530, 
    9209, 9531, 9774, 9854, 9759, 10113, 9930, 9930, 10018, 9801, 9646, 9701, 
    9769, 9879, 9739, 9625, 9862, 10046, 9930, 9930, 9930, 9930, 9930, 9930, 
    9930, 9930,
  9674, 9395, 8987, 9118, 8629, 8204, 8318, 8578, 8822, 8972, 8822, 8492, 
    8789, 8954, 9000, 8345, 8086, 8855, 9506, 8915, 8756, 8748, 9284, 9587, 
    9776, 9822, 9939, 10018, 10018, 10018, 10018, 10018, 9986, 9943, 9932, 
    9931, 9951, 9860, 9840, 9943, 9971, 9980, 9939, 9834, 9854, 9860, 9936, 
    9870, 9884, 9861, 9999, 9810, 9632, 9912, 9992, 10015, 10018, 10018, 
    10018, 10018, 9905, 9830, 9708, 9810, 9888, 9729, 9487, 9403, 9600, 9306, 
    9642, 9645, 9804, 9976, 9884, 10105, 9930, 9930, 9987, 9774, 9580, 9859, 
    9861, 9932, 9897, 9849, 10046, 9930, 9930, 9930, 9930, 9930, 9930, 9930, 
    9930, 9930,
  9796, 9395, 9154, 8790, 8781, 8452, 8416, 8609, 8831, 9004, 8977, 8785, 
    8709, 8783, 8988, 8720, 8227, 7646, 9474, 9049, 8770, 8968, 9273, 9510, 
    9814, 9960, 9992, 10018, 10018, 10018, 9990, 10018, 10018, 10018, 9957, 
    10018, 9977, 9973, 9854, 9923, 9999, 10008, 9994, 10008, 9969, 9980, 
    9992, 9854, 9954, 9971, 9964, 9900, 9893, 9906, 10018, 10018, 10018, 
    10018, 10018, 10018, 9668, 9625, 9746, 9814, 9884, 9849, 9349, 9149, 
    9587, 9447, 9862, 9862, 9939, 10069, 10084, 9930, 9930, 9930, 9979, 9780, 
    9783, 9860, 9909, 9918, 10020, 10053, 9930, 9930, 9930, 9930, 9930, 9930, 
    9930, 9930, 9930, 9930,
  9796, 9701, 9519, 9040, 8709, 8382, 8376, 8565, 8631, 8767, 8935, 8693, 
    8967, 8620, 8450, 8842, 8314, 8427, 9306, 9066, 8801, 8989, 9439, 9575, 
    9870, 9974, 10018, 10018, 10018, 10018, 10010, 10018, 10018, 10018, 
    10018, 10018, 10018, 10008, 10002, 9971, 10018, 10018, 10010, 10018, 
    10018, 10018, 9987, 9948, 10010, 10008, 10008, 10018, 9971, 10002, 10018, 
    10018, 10018, 10018, 10018, 10018, 9948, 9756, 9736, 9767, 9838, 9646, 
    9607, 9371, 9382, 9688, 9977, 10013, 10036, 10051, 10084, 9930, 9930, 
    10121, 9879, 9693, 9711, 10008, 10043, 9882, 10020, 10084, 9930, 9930, 
    9930, 9930, 9930, 9930, 9930, 9930, 9930, 9930,
  9776, 9824, 9621, 9177, 8977, 8519, 8424, 8464, 8881, 8987, 9030, 8938, 
    8680, 8675, 8480, 8770, 8548, 8927, 9306, 9215, 8510, 9028, 9258, 9762, 
    9986, 10004, 10018, 10018, 10018, 10018, 10018, 10018, 10018, 10018, 
    10018, 10018, 10010, 10018, 10018, 10010, 10018, 10018, 10018, 10018, 
    10018, 10018, 10018, 10015, 10014, 10018, 10018, 10018, 10018, 10018, 
    10018, 10018, 10018, 10018, 10018, 10102, 10009, 9854, 9646, 9592, 9731, 
    9547, 9601, 9681, 9649, 9751, 10041, 10080, 10051, 10036, 10111, 10102, 
    9930, 9930, 9943, 9514, 9711, 10084, 10084, 10084, 9930, 9930, 9930, 
    9930, 9930, 9930, 9930, 9930, 9930, 9930, 9930, 9930,
  9796, 9804, 9796, 9485, 9008, 8709, 8356, 8533, 8912, 8808, 8876, 8740, 
    8658, 8852, 8658, 8896, 8989, 9145, 9245, 8667, 8401, 9313, 9462, 9872, 
    9964, 10018, 10018, 10018, 10018, 10018, 10018, 10018, 10018, 10018, 
    10018, 10018, 9997, 10018, 10018, 10018, 10018, 10018, 10018, 10018, 
    10018, 10018, 10018, 10018, 10018, 10018, 10018, 10018, 10018, 10018, 
    10018, 10018, 10018, 10018, 10018, 10018, 10007, 9704, 9625, 9447, 9729, 
    9620, 9563, 9894, 9931, 9837, 10029, 10084, 10084, 10076, 10064, 10064, 
    10126, 10084, 9715, 9546, 9923, 10084, 9930, 9930, 9930, 9930, 9930, 
    9930, 9930, 9930, 9930, 9930, 9930, 9930, 9930, 9930,
  9796, 9813, 9826, 9612, 9145, 8740, 8378, 8508, 8750, 8770, 8724, 8651, 
    8598, 9316, 8466, 8903, 9072, 9200, 9397, 8759, 8876, 8927, 9694, 9974, 
    10007, 10018, 10018, 9942, 9928, 10018, 9983, 10018, 10018, 10018, 10018, 
    10018, 10018, 10002, 10018, 10018, 10018, 10018, 10018, 10018, 10018, 
    10018, 10018, 10018, 10018, 10018, 10018, 10018, 10018, 10018, 10018, 
    10018, 10018, 10018, 10046, 10130, 10130, 9970, 9614, 9546, 9852, 9687, 
    9731, 9838, 10095, 10085, 10084, 9930, 9930, 10084, 10097, 10101, 10084, 
    10084, 10074, 10084, 10084, 9930, 9930, 9930, 9930, 9930, 9930, 9930, 
    9930, 9930, 9930, 9930, 9930, 9930, 9930, 9930,
  9796, 9832, 9832, 9712, 9156, 8699, 8423, 8568, 8803, 8772, 8819, 8159, 
    8829, 8791, 8629, 9134, 9142, 9494, 9201, 8559, 8770, 9349, 9837, 9870, 
    10018, 9941, 9963, 9847, 9847, 9951, 9969, 10009, 10018, 10018, 10018, 
    10018, 10018, 10004, 10018, 10012, 10018, 10018, 10018, 10018, 10018, 
    10018, 10018, 10018, 10018, 10018, 10018, 10018, 10018, 10018, 10018, 
    10018, 10018, 10046, 10054, 10054, 10074, 10029, 9882, 9817, 9838, 9764, 
    9979, 10067, 10084, 10084, 9930, 9930, 9930, 10084, 10084, 10084, 10084, 
    10084, 10084, 10084, 10084, 10084, 9930, 9930, 9930, 9930, 9930, 9930, 
    9930, 9930, 9930, 9930, 9930, 9930, 9930, 9930,
  9796, 9832, 9832, 9792, 9177, 8815, 8682, 8548, 8827, 8904, 8678, 8318, 
    8663, 9023, 8977, 9049, 9109, 9448, 8915, 8658, 8924, 9662, 9936, 9990, 
    10018, 9969, 9790, 9822, 9897, 9943, 9971, 9960, 10012, 10018, 10018, 
    10018, 10018, 10018, 10018, 9990, 10018, 10018, 10018, 10018, 10018, 
    10018, 10018, 10018, 10018, 10018, 10018, 10018, 10018, 10018, 10018, 
    10018, 10018, 10046, 10054, 10054, 10116, 10121, 10084, 9985, 10025, 
    10084, 10084, 10084, 10084, 10084, 10084, 10084, 10084, 10084, 10084, 
    10084, 10084, 10084, 10084, 10084, 10084, 10084, 10084, 9930, 9930, 9930, 
    9930, 9930, 10130, 10130, 9930, 9930, 9930, 9930, 9930, 9930,
  9796, 9832, 9832, 9806, 9220, 8781, 8700, 8691, 8770, 8702, 8729, 8440, 
    8585, 9019, 8852, 9395, 9399, 9316, 8482, 8372, 9135, 9701, 9883, 10015, 
    9907, 9907, 9627, 9748, 9799, 9894, 9951, 9980, 9974, 10015, 10018, 
    10018, 10018, 10018, 10018, 10010, 10018, 10018, 10018, 10018, 10018, 
    10018, 10018, 10018, 10018, 10018, 10018, 10018, 10018, 10018, 10018, 
    10018, 10018, 10018, 10054, 10092, 10121, 10084, 10084, 10084, 9930, 
    9930, 10084, 10084, 10084, 10084, 10084, 10084, 10084, 9930, 9930, 10084, 
    10084, 10084, 10084, 10084, 10084, 10084, 9930, 9930, 9930, 9930, 9930, 
    10130, 10092, 10130, 9930, 10084, 9930, 9930, 9930, 9930,
  9796, 9832, 9832, 9636, 9093, 8663, 8742, 8858, 8874, 8629, 8494, 8275, 
    8739, 8683, 9060, 9614, 9749, 9487, 8645, 8631, 9313, 9558, 9946, 10018, 
    9920, 9849, 9580, 9734, 9801, 9743, 9932, 9980, 9980, 10008, 10018, 
    10018, 10018, 10018, 10018, 10018, 10018, 10018, 10018, 10018, 10018, 
    10018, 10018, 10018, 10018, 10018, 10018, 10018, 10018, 10018, 10018, 
    10018, 10018, 10018, 10046, 10092, 10084, 10084, 10084, 10084, 10084, 
    10084, 10084, 10084, 10084, 10084, 10084, 10084, 10084, 10084, 10084, 
    10084, 10084, 10084, 10084, 10084, 10084, 10084, 10084, 10084, 9930, 
    9930, 9930, 9930, 9946, 9906, 9879, 10084, 10084, 9930, 9930, 9930,
  9796, 9824, 9832, 9317, 9082, 9213, 8809, 8795, 8852, 8856, 8471, 8415, 
    8548, 8711, 8740, 9511, 9794, 8991, 8490, 8559, 9448, 9731, 9981, 10018, 
    10018, 9858, 9616, 9601, 9721, 9724, 9890, 9936, 10008, 10015, 10018, 
    10018, 10018, 10018, 10018, 10018, 10018, 10018, 10018, 10018, 10018, 
    10018, 10018, 10018, 10018, 10018, 10018, 10018, 10018, 10018, 10018, 
    10018, 10018, 10018, 10090, 9930, 9930, 10084, 10084, 10084, 10084, 
    10084, 10084, 10084, 10084, 10084, 10084, 10084, 10084, 10084, 10084, 
    10084, 10084, 10084, 10084, 10084, 10084, 10084, 10084, 10084, 10084, 
    9930, 9930, 9930, 10084, 9832, 9796, 9930, 10084, 9930, 9930, 9930 ;

 TPW =
  121, 119, 83, 108, 89, 78, 81, 84, 96, 95, 93, 108, 98, 110, 109, 91, 85, 
    119, 144, 145, 150, 155, 200, 256, 305, 318, 317, 328, 347, 348, 339, 
    335, 260, 342, 344, 337, 328, 321, 302, 316, 310, 257, 259, 197, 229, 
    257, 238, 253, 253, 247, 209, 174, 231, 265, 298, 281, 195, 198, 220, 
    270, 224, 211, 202, 225, 184, 183, 184, 164, 155, 145, 133, 181, 153, 
    124, 140, 120, 85, 81, 118, 104, 115, 126, 134, 132, 105, 115, 113, 105, 
    115, 115, 111, 100, 107, 126, 118, 142,
  126, 104, 90, 106, 77, 68, 73, 85, 85, 95, 91, 92, 90, 91, 97, 89, 93, 118, 
    180, 161, 169, 221, 237, 296, 313, 333, 319, 346, 323, 328, 352, 340, 
    335, 329, 331, 338, 341, 313, 314, 335, 349, 280, 143, 202, 270, 263, 
    333, 343, 306, 271, 223, 219, 293, 280, 283, 257, 150, 179, 202, 240, 
    222, 206, 190, 184, 184, 156, 149, 144, 133, 120, 129, 129, 120, 141, 
    124, 108, 86, 85, 119, 130, 110, 118, 119, 119, 144, 116, 109, 93, 107, 
    104, 108, 96, 103, 110, 101, 92,
  122, 108, 95, 87, 82, 70, 71, 73, 90, 98, 99, 90, 81, 88, 101, 111, 109, 
    122, 193, 194, 184, 252, 294, 311, 341, 372, 349, 334, 304, 313, 338, 
    340, 340, 329, 320, 298, 311, 289, 259, 245, 250, 209, 135, 218, 230, 
    225, 242, 230, 347, 258, 301, 301, 276, 300, 227, 204, 188, 157, 175, 
    214, 190, 192, 167, 166, 137, 157, 146, 132, 136, 130, 143, 124, 125, 
    129, 104, 80, 80, 75, 126, 138, 134, 152, 143, 140, 144, 116, 91, 112, 
    106, 104, 113, 120, 106, 105, 95, 95,
  128, 123, 123, 100, 91, 73, 79, 76, 82, 91, 90, 81, 96, 84, 104, 142, 159, 
    177, 224, 230, 265, 262, 314, 312, 354, 349, 355, 320, 316, 337, 335, 
    361, 343, 323, 296, 294, 256, 261, 265, 174, 195, 154, 136, 120, 198, 
    164, 172, 213, 142, 182, 262, 278, 245, 211, 188, 184, 182, 166, 158, 
    201, 167, 165, 155, 143, 130, 123, 130, 116, 128, 125, 127, 128, 126, 
    119, 90, 81, 87, 109, 126, 135, 153, 150, 135, 109, 108, 103, 89, 105, 
    107, 111, 110, 118, 106, 105, 96, 85,
  129, 121, 127, 111, 99, 77, 69, 77, 86, 88, 88, 95, 97, 107, 119, 218, 250, 
    280, 329, 308, 240, 280, 281, 345, 358, 337, 323, 311, 306, 295, 314, 
    309, 285, 270, 273, 289, 257, 226, 228, 227, 140, 145, 194, 202, 187, 
    169, 194, 202, 217, 217, 210, 252, 201, 194, 183, 158, 158, 199, 182, 
    148, 159, 160, 139, 130, 145, 120, 141, 127, 125, 133, 142, 123, 120, 
    112, 94, 115, 80, 80, 126, 125, 137, 119, 101, 101, 88, 88, 95, 111, 112, 
    116, 117, 112, 129, 117, 94, 119,
  119, 129, 132, 125, 102, 92, 69, 82, 87, 85, 92, 87, 107, 134, 175, 282, 
    293, 282, 339, 261, 221, 299, 314, 350, 325, 320, 308, 321, 315, 308, 
    324, 296, 268, 253, 243, 255, 251, 235, 225, 212, 225, 148, 192, 176, 
    113, 182, 201, 216, 214, 214, 233, 214, 187, 195, 191, 160, 168, 177, 
    160, 163, 149, 153, 134, 117, 146, 126, 130, 124, 139, 140, 128, 103, 99, 
    96, 95, 122, 115, 89, 127, 140, 116, 99, 84, 82, 88, 96, 111, 106, 106, 
    105, 108, 116, 123, 122, 116, 123,
  119, 122, 131, 144, 115, 83, 72, 79, 81, 88, 103, 105, 114, 189, 210, 261, 
    287, 339, 337, 248, 258, 273, 341, 365, 328, 305, 305, 323, 312, 310, 
    337, 318, 308, 280, 254, 248, 244, 253, 304, 163, 124, 198, 182, 182, 
    184, 192, 195, 202, 211, 191, 192, 211, 192, 174, 157, 187, 151, 153, 
    149, 146, 142, 143, 126, 132, 143, 129, 104, 118, 110, 107, 99, 80, 85, 
    91, 120, 120, 97, 98, 115, 102, 98, 78, 87, 88, 96, 112, 120, 115, 107, 
    103, 114, 118, 118, 118, 113, 120,
  121, 127, 134, 141, 109, 90, 77, 82, 84, 96, 129, 103, 141, 232, 245, 273, 
    278, 337, 274, 229, 244, 299, 331, 324, 317, 315, 319, 303, 279, 299, 
    324, 313, 313, 293, 263, 266, 254, 246, 257, 236, 229, 225, 188, 192, 
    191, 197, 194, 187, 189, 185, 205, 186, 188, 169, 179, 174, 148, 152, 
    137, 144, 137, 127, 119, 126, 115, 101, 118, 120, 94, 98, 86, 85, 75, 96, 
    95, 98, 100, 105, 106, 102, 105, 107, 113, 86, 110, 108, 122, 113, 110, 
    96, 108, 120, 130, 121, 123, 113,
  126, 125, 116, 114, 106, 92, 87, 77, 89, 106, 122, 145, 198, 294, 277, 264, 
    267, 258, 263, 229, 257, 303, 322, 327, 341, 316, 284, 285, 270, 280, 
    283, 287, 265, 271, 268, 237, 235, 230, 252, 270, 244, 277, 190, 195, 
    185, 188, 184, 195, 192, 191, 195, 201, 188, 172, 142, 140, 147, 135, 
    128, 147, 143, 140, 130, 141, 116, 110, 90, 91, 94, 89, 94, 98, 99, 100, 
    95, 93, 98, 103, 110, 106, 106, 107, 103, 102, 98, 112, 120, 118, 107, 
    107, 107, 114, 126, 130, 119, 120,
  117, 131, 120, 119, 103, 82, 87, 94, 124, 122, 182, 189, 243, 286, 265, 
    276, 269, 286, 213, 204, 264, 326, 329, 323, 314, 327, 308, 281, 267, 
    262, 281, 277, 246, 235, 242, 248, 240, 222, 246, 251, 237, 239, 184, 
    183, 200, 195, 128, 194, 193, 196, 201, 191, 186, 162, 144, 145, 145, 
    138, 129, 135, 142, 130, 118, 104, 97, 91, 102, 98, 97, 99, 97, 99, 101, 
    83, 84, 97, 100, 103, 104, 99, 106, 105, 103, 92, 94, 106, 103, 109, 119, 
    116, 128, 95, 133, 126, 124, 125,
  114, 117, 126, 116, 89, 83, 93, 117, 144, 144, 198, 214, 275, 240, 207, 
    267, 319, 309, 217, 207, 281, 301, 343, 318, 321, 297, 278, 250, 254, 
    180, 244, 245, 231, 231, 210, 232, 226, 256, 227, 223, 219, 217, 190, 
    204, 160, 188, 188, 189, 199, 185, 169, 187, 177, 145, 179, 156, 135, 
    128, 132, 135, 120, 126, 116, 111, 105, 103, 99, 101, 102, 97, 89, 90, 
    92, 92, 96, 95, 96, 107, 100, 102, 104, 103, 98, 97, 116, 100, 112, 101, 
    115, 116, 111, 113, 103, 122, 125, 120,
  107, 127, 140, 108, 98, 102, 118, 140, 185, 249, 221, 164, 224, 227, 192, 
    359, 315, 269, 206, 187, 247, 277, 300, 291, 305, 287, 254, 251, 247, 
    252, 258, 241, 235, 259, 249, 270, 208, 233, 220, 230, 218, 215, 207, 
    196, 185, 166, 151, 178, 188, 198, 171, 186, 151, 164, 166, 168, 127, 
    123, 122, 112, 102, 125, 121, 106, 103, 102, 102, 100, 98, 96, 91, 88, 
    92, 95, 96, 96, 98, 99, 100, 100, 101, 106, 111, 106, 103, 113, 126, 121, 
    110, 118, 124, 139, 95, 127, 130, 113 ;

 TSkin =
  31080, 31174, 30955, 30845, 30819, 30888, 30927, 31227, 31114, 31041, 
    30909, 30487, 30539, 30649, 30279, 30465, 30360, 30331, 30192, 30316, 
    30332, 30342, 30004, 29642, 29549, 29674, 29268, 29132, 28826, 28993, 
    29216, 29406, 29371, 29443, 29299, 29231, 29103, 28753, 28811, 28783, 
    28596, 28227, 28031, 28044, 28174, 28175, 27934, 28100, 28156, 28319, 
    27863, 28415, 28535, 28601, 28725, 28732, 28765, 28327, 28359, 28732, 
    28960, 28950, 29035, 29053, 28884, 29008, 29053, 29049, 29029, 28755, 
    28822, 28376, 28665, 28775, 28576, 27286, 26589, 26723, 27882, 28906, 
    28851, 28713, 28784, 28611, 28873, 28675, 28232, 27503, 27425, 27538, 
    27878, 27820, 27750, 27842, 27630, 28100,
  31057, 31233, 31072, 30822, 30979, 30690, 30837, 30842, 30914, 31022, 
    30942, 30578, 30645, 30599, 30348, 30418, 30148, 30059, 29915, 30257, 
    30150, 30088, 29617, 29306, 29240, 29462, 29282, 28951, 28563, 28738, 
    28949, 28991, 28824, 28839, 29223, 28931, 29013, 28675, 28864, 28960, 
    28772, 27989, 28036, 29110, 28387, 28350, 28919, 29013, 28604, 28440, 
    29456, 29621, 28772, 28720, 28793, 28453, 28290, 27958, 27950, 28728, 
    29015, 29174, 29054, 29118, 28949, 29108, 29147, 29341, 28945, 28839, 
    28745, 28622, 28709, 28497, 28062, 26834, 26566, 27139, 28258, 28896, 
    28855, 28625, 28562, 28588, 28458, 28234, 27460, 27431, 27593, 27585, 
    27982, 27848, 27901, 27975, 27718, 27320,
  31165, 31176, 31106, 30857, 30777, 30668, 30808, 30789, 30855, 30974, 
    30797, 30698, 30554, 30552, 30218, 30292, 30339, 29964, 30120, 30283, 
    30182, 29796, 29403, 29226, 29157, 29265, 29093, 28612, 28925, 29249, 
    29626, 29572, 29475, 29275, 29002, 28961, 28799, 28596, 28582, 29580, 
    29338, 27898, 28121, 28993, 29022, 29266, 29409, 29499, 28673, 29419, 
    29411, 29438, 29489, 29189, 29126, 28900, 28514, 27737, 27853, 28359, 
    28968, 29116, 29089, 29037, 28914, 28986, 29195, 29089, 29101, 28981, 
    28828, 28819, 28567, 27966, 28297, 26990, 26709, 26918, 28268, 29124, 
    28976, 28555, 28344, 28297, 27686, 27191, 27006, 27116, 27634, 27723, 
    27885, 27960, 27918, 27719, 27835, 27466,
  31212, 31286, 31062, 31049, 30911, 30574, 30803, 30666, 30865, 30976, 
    30853, 30967, 30555, 30396, 30318, 30259, 30069, 30102, 29934, 30112, 
    29955, 29693, 29353, 29160, 29256, 28986, 28840, 28783, 28889, 29374, 
    29787, 30194, 29443, 28898, 28866, 28523, 28472, 28048, 28048, 28318, 
    28188, 27968, 28186, 27979, 28623, 27971, 28037, 28712, 28116, 28283, 
    28757, 29206, 29022, 28764, 28650, 28415, 28232, 27684, 27774, 28045, 
    28576, 28959, 29116, 29067, 29092, 29084, 29100, 29018, 28765, 28779, 
    28745, 28682, 28402, 27730, 28172, 26866, 26666, 26699, 28467, 29406, 
    28877, 28031, 27366, 27822, 27125, 27912, 27122, 27222, 27666, 27817, 
    27847, 28078, 27840, 27673, 27733, 27739,
  31299, 31060, 31153, 31024, 30710, 30679, 30749, 30803, 30814, 30991, 
    30623, 30740, 30649, 30516, 30360, 30035, 29825, 29977, 30225, 29992, 
    29575, 29494, 29300, 29226, 29240, 28805, 28910, 29203, 29283, 29598, 
    29331, 29116, 28753, 28419, 28462, 28482, 28417, 28236, 28178, 29050, 
    27966, 27821, 28730, 28680, 27514, 27938, 27577, 28636, 28719, 27856, 
    28153, 28028, 28548, 28295, 28218, 27858, 27552, 27521, 27583, 27745, 
    28285, 29020, 28950, 29160, 28854, 28945, 28701, 28708, 28861, 28946, 
    28606, 27784, 27508, 27394, 27254, 27083, 26971, 27384, 28201, 29203, 
    28079, 28169, 28101, 27916, 26842, 26859, 27240, 27357, 27614, 27814, 
    27820, 28024, 28235, 28218, 27843, 28570,
  31363, 31308, 31263, 31040, 30821, 30844, 30636, 30637, 30778, 30703, 
    30708, 30755, 30741, 30161, 30156, 29760, 29752, 30629, 30567, 29815, 
    29699, 29481, 29269, 29132, 29023, 28845, 29008, 29285, 29287, 29161, 
    28986, 28873, 29590, 29488, 29441, 29398, 29403, 29094, 29060, 29048, 
    28582, 27979, 28558, 28520, 27898, 27749, 28532, 28725, 28105, 28787, 
    28806, 28606, 27806, 28319, 28114, 27485, 27484, 27238, 27529, 27698, 
    28047, 28871, 29151, 28916, 28772, 28891, 28924, 28685, 28856, 28351, 
    27001, 28170, 28162, 27116, 27466, 28142, 26878, 28261, 27535, 28356, 
    26785, 27988, 26971, 26936, 26950, 27141, 27385, 27607, 27513, 27629, 
    27718, 28055, 28090, 28121, 28389, 28577,
  31360, 31327, 31102, 30879, 30694, 30907, 30730, 30766, 30642, 30739, 
    30774, 30674, 30569, 30066, 30138, 29733, 29257, 30408, 29919, 29834, 
    29738, 29694, 29498, 29188, 28728, 28815, 29239, 29065, 28830, 28649, 
    28857, 29292, 29539, 29466, 29347, 29339, 29260, 29351, 28565, 28308, 
    28199, 28792, 28704, 28426, 28404, 28476, 28462, 28491, 28404, 28036, 
    27990, 27651, 27924, 27833, 27393, 27449, 27277, 27078, 27398, 27512, 
    27880, 28498, 28844, 28913, 29041, 28758, 28860, 28346, 27293, 26772, 
    28138, 26734, 26570, 28253, 27315, 27779, 28341, 28142, 27204, 28325, 
    28129, 26701, 26758, 26944, 27371, 27524, 27639, 27688, 27434, 27608, 
    27709, 28050, 28103, 28234, 28253, 28418,
  31431, 31279, 31212, 31146, 30835, 30944, 30875, 30722, 30640, 30675, 
    30762, 30714, 30457, 30007, 29501, 29310, 29255, 29726, 29611, 30017, 
    29867, 29685, 29357, 29171, 28732, 28811, 28771, 28631, 28626, 28621, 
    28520, 28595, 28816, 29034, 28851, 28781, 29188, 29228, 28513, 28342, 
    28338, 28229, 28666, 28399, 28263, 28470, 28340, 28217, 28220, 28299, 
    28335, 28159, 28040, 27720, 27343, 26986, 27186, 27160, 27279, 27344, 
    27567, 28050, 28621, 28761, 28665, 28720, 28133, 26862, 28048, 28066, 
    26409, 26384, 26780, 28152, 28289, 28324, 28294, 28153, 28123, 28093, 
    28113, 28080, 27961, 27250, 27643, 27907, 27715, 27749, 27420, 27608, 
    27685, 28094, 27993, 28133, 28310, 28424,
  31468, 31330, 31303, 31147, 30970, 30816, 30965, 30887, 30710, 30405, 
    30383, 30223, 30080, 29682, 29372, 29521, 29564, 29462, 29446, 29473, 
    29188, 29395, 29829, 29057, 28765, 28649, 28904, 28678, 28562, 28611, 
    28474, 28224, 28414, 28051, 28394, 28159, 28232, 28408, 28235, 28559, 
    28219, 27907, 28077, 28274, 28230, 28347, 28365, 28117, 28144, 28134, 
    28195, 27683, 28039, 28017, 27154, 27049, 27191, 27190, 27105, 27196, 
    27179, 27243, 28597, 27139, 26942, 28413, 28177, 28205, 28001, 28224, 
    28167, 28156, 28260, 28166, 28210, 28152, 28349, 28252, 28161, 28212, 
    28143, 28121, 27980, 27725, 27780, 27551, 27553, 27366, 27223, 27502, 
    27822, 28078, 28046, 27943, 28036, 28298,
  31516, 31177, 31268, 31049, 30889, 30765, 30876, 30809, 30796, 30438, 
    30181, 30151, 29749, 29044, 29627, 30051, 29983, 29367, 29444, 29265, 
    29153, 29155, 29004, 28864, 28722, 28914, 28897, 28808, 28504, 28592, 
    28453, 28406, 28299, 28203, 27986, 28182, 28218, 28927, 28749, 28357, 
    28282, 27873, 27822, 27412, 28091, 28110, 27905, 28254, 28202, 28327, 
    27903, 28014, 28421, 27773, 27446, 27443, 27628, 27226, 27172, 27181, 
    26790, 28389, 28290, 28294, 26009, 26524, 28093, 28072, 28208, 28187, 
    28155, 28092, 28197, 26497, 26421, 28106, 28157, 28205, 28137, 28072, 
    28108, 28035, 27821, 27825, 27749, 27502, 27460, 27061, 27463, 27743, 
    27945, 27764, 27978, 27967, 27967, 28221,
  31617, 31425, 31230, 30996, 30933, 30673, 30753, 30725, 30613, 30508, 
    29999, 29598, 29667, 29230, 29745, 29756, 29954, 29421, 29374, 29379, 
    29071, 29065, 29014, 28954, 28962, 28921, 28713, 28527, 28579, 28191, 
    28374, 28330, 28310, 27725, 27810, 27947, 28830, 28379, 28358, 28163, 
    27931, 27774, 27922, 27882, 27738, 28105, 28207, 28286, 28301, 28047, 
    28101, 28431, 28389, 27689, 27589, 27654, 27696, 27405, 27278, 26441, 
    28399, 28379, 28220, 28191, 28242, 28217, 28132, 28177, 28066, 28134, 
    28172, 28161, 28119, 28088, 28123, 28092, 28105, 28108, 28200, 28088, 
    28035, 28060, 28022, 27908, 27335, 27444, 27217, 27137, 27523, 28359, 
    28235, 27851, 27695, 27843, 28055, 28128,
  31457, 31285, 31015, 31124, 30935, 31012, 30715, 30574, 30224, 29910, 
    29416, 29904, 29853, 29899, 30006, 29934, 29950, 29375, 29102, 29211, 
    29018, 28945, 28722, 28727, 28955, 28818, 28819, 28744, 28559, 28393, 
    28099, 28354, 28367, 28052, 28089, 27822, 28715, 27813, 27726, 27676, 
    27754, 27655, 27725, 27658, 27781, 27607, 27495, 28271, 28307, 28580, 
    28018, 28172, 27723, 27818, 27886, 27616, 27766, 27559, 26846, 26741, 
    26674, 28436, 28212, 28249, 28199, 28117, 28061, 28133, 28014, 28171, 
    28087, 28121, 28025, 28027, 28105, 28037, 27963, 28024, 28101, 28077, 
    27967, 27996, 27954, 27960, 27824, 27331, 27305, 27211, 27795, 28335, 
    28165, 27753, 27668, 27753, 28025, 27358 ;

 WindDir =
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888 ;

 WindSp =
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888 ;

 WindU =
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888 ;

 WindV =
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, 
    -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888, -888 ;

 YM =
  28616, 28565, 27757, 26985, 25698, 24124, 22683, 22188, 22092, 22443, 
    22808, 23615, 24611, 25870, 26382, 28476, 28644, 27831, 27278, 26697, 
    25900, 25117,
  28582, 28533, 27831, 27057, 25869, 24263, 22769, 22211, 22092, 22492, 
    22782, 23574, 24719, 25684, 26438, 28521, 28718, 27788, 27250, 26747, 
    25888, 24963,
  28495, 28463, 27740, 27138, 25972, 24350, 22901, 22279, 22124, 22448, 
    22862, 23566, 24465, 25690, 26834, 28429, 28532, 27795, 27188, 26703, 
    25913, 24963,
  28393, 28393, 27754, 27154, 26043, 24462, 22914, 22282, 22091, 22480, 
    22853, 23507, 24472, 25690, 26532, 28303, 28488, 27679, 27132, 26585, 
    25893, 24942,
  28314, 28346, 27717, 27195, 26132, 24571, 23011, 22267, 22129, 22508, 
    22878, 23467, 24401, 25710, 26454, 28262, 28426, 27651, 27035, 26448, 
    25701, 24869,
  28286, 28333, 27742, 27210, 26220, 24663, 23060, 22387, 22170, 22462, 
    22810, 23497, 24529, 25583, 26626, 28245, 28395, 27607, 27029, 26373, 
    25556, 24721,
  28326, 28368, 27804, 27319, 26315, 24800, 23129, 22386, 22137, 22439, 
    22824, 23459, 24412, 25485, 26391, 28460, 28544, 27723, 27001, 26373, 
    25511, 24627,
  28411, 28441, 28018, 27459, 26469, 24840, 23188, 22433, 22160, 22447, 
    22815, 23481, 24420, 25610, 26292, 28566, 28756, 27766, 27070, 26317, 
    25447, 24634,
  28488, 28508, 28079, 27560, 26532, 24951, 23274, 22480, 22151, 22407, 
    22818, 23420, 24417, 25513, 26432, 28642, 28762, 27707, 27001, 26373, 
    25389, 24486,
  28506, 28524, 28140, 27609, 26585, 24999, 23347, 22518, 22189, 22415, 
    22820, 23448, 24424, 25482, 26479, 28628, 28687, 27701, 26910, 26217, 
    25185, 24238,
  28461, 28485, 28072, 27598, 26579, 25043, 23392, 22559, 22189, 22389, 
    22754, 23447, 24355, 25422, 26376, 28582, 28706, 27521, 26779, 25987, 
    24937, 24137,
  28387, 28416, 27940, 27496, 26531, 25037, 23423, 22580, 22191, 22397, 
    22942, 23384, 24355, 25410, 26420, 28410, 28388, 27354, 26642, 25757, 
    24880, 24004,
  28303, 28325, 27856, 27485, 26592, 25155, 23481, 22630, 22217, 22445, 
    22862, 23381, 24300, 25293, 26591, 28217, 28214, 27354, 26545, 25738, 
    24688, 23970,
  28199, 28208, 27899, 27488, 26640, 25189, 23513, 22641, 22261, 22494, 
    22842, 23431, 24549, 25533, 26085, 28251, 28388, 27441, 26662, 25831, 
    24784, 24016,
  28072, 28078, 27832, 27469, 26642, 25250, 23610, 22673, 22225, 22396, 
    22907, 23370, 24302, 25519, 26438, 28223, 28376, 27499, 26731, 25943, 
    24841, 24036,
  27954, 27973, 27721, 27407, 26628, 25275, 23596, 22714, 22281, 22442, 
    22776, 23367, 24290, 25360, 26610, 28032, 28264, 27549, 26821, 25935, 
    25000, 24216,
  27883, 27916, 27625, 27269, 26639, 25261, 23651, 22758, 22307, 22467, 
    22812, 23435, 24211, 25437, 26559, 27876, 28190, 27441, 26641, 25804, 
    24859, 24196,
  27867, 27905, 27567, 27321, 26663, 25340, 23692, 22749, 22289, 22430, 
    22806, 23448, 24146, 25453, 26376, 27869, 28207, 27253, 26434, 25613, 
    24821, 24109,
  27887, 27926, 27688, 27409, 26714, 25384, 23755, 22790, 22303, 22429, 
    22761, 23318, 24358, 25167, 26259, 27985, 28220, 27123, 26324, 25594, 
    24795, 24216,
  27919, 27970, 27749, 27439, 26754, 25423, 23772, 22840, 22362, 22394, 
    22829, 23323, 24185, 25418, 26467, 28034, 28046, 26870, 26088, 25420, 
    24807, 24275,
  27951, 28024, 27826, 27476, 26785, 25465, 23796, 22831, 22332, 22460, 
    22723, 23310, 24353, 25425, 26585, 28051, 28026, 26819, 26096, 25345, 
    24654, 24074,
  27988, 28073, 27812, 27496, 26788, 25493, 23813, 22863, 22396, 22457, 
    22780, 23348, 24281, 25308, 26551, 28140, 28089, 26812, 26019, 25319, 
    24718, 24087,
  28025, 28096, 27764, 27428, 26771, 25496, 23858, 22928, 22361, 22391, 
    22765, 23333, 24165, 25299, 26341, 28084, 27965, 26740, 26040, 25388, 
    24685, 24094,
  28017, 28040, 27693, 27423, 26731, 25484, 23865, 22921, 22405, 22379, 
    22810, 23360, 24327, 25399, 26638, 27970, 27741, 26675, 26101, 25469, 
    24768, 24221,
  27886, 27839, 27735, 27401, 26699, 25501, 23906, 22912, 22431, 22442, 
    22713, 23230, 24186, 25317, 26432, 28037, 27741, 26638, 26046, 25449, 
    24736, 24200,
  27606, 27482, 27690, 27350, 26734, 25518, 23910, 22960, 22422, 22390, 
    22722, 23266, 24119, 25110, 26319, 28026, 27753, 26559, 25943, 25424, 
    24768, 24080,
  27247, 27074, 27368, 27218, 26659, 25481, 23941, 22956, 22442, 22419, 
    22822, 23334, 24156, 25457, 26191, 27735, 27629, 26566, 25922, 25368, 
    24665, 24160,
  26957, 26771, 27041, 27001, 26585, 25442, 23944, 22986, 22430, 22427, 
    22616, 23240, 24203, 25317, 25973, 27399, 27591, 26501, 25935, 25412, 
    24704, 24179,
  26862, 26676, 26825, 26868, 26541, 25470, 23958, 23000, 22438, 22467, 
    22741, 23291, 24119, 25249, 26226, 27248, 27398, 26443, 25922, 25399, 
    24678, 24065,
  26984, 26795, 27023, 27016, 26573, 25537, 23975, 22985, 22506, 22478, 
    22744, 23270, 23958, 25466, 26284, 27363, 27442, 26428, 25879, 25361, 
    24639, 24079,
  27229, 27055, 27312, 27185, 26662, 25537, 24006, 23050, 22502, 22490, 
    22824, 23326, 24227, 25189, 26326, 27632, 27604, 26485, 25866, 25374, 
    24652, 24105,
  27463, 27343, 27403, 27274, 26725, 25559, 23995, 23064, 22482, 22470, 
    22752, 23290, 24111, 25158, 26531, 27806, 27660, 26443, 25825, 25230, 
    24658, 24145,
  27613, 27553, 27449, 27296, 26713, 25581, 24023, 23041, 22531, 22481, 
    22755, 23358, 24237, 25342, 26345, 27809, 27734, 26370, 25810, 25230, 
    24677, 24098,
  27682, 27640, 27594, 27376, 26760, 25601, 24065, 23055, 22555, 22526, 
    22737, 23330, 24081, 25300, 26371, 27842, 27616, 26370, 25824, 25280, 
    24600, 24085,
  27701, 27640, 27679, 27371, 26742, 25576, 24027, 23058, 22534, 22546, 
    22791, 23376, 24163, 25316, 26299, 27956, 27504, 26363, 25817, 25212, 
    24575, 24124,
  27686, 27614, 27698, 27368, 26784, 25545, 24033, 23090, 22528, 22492, 
    22817, 23350, 24110, 25255, 26306, 27912, 27466, 26370, 25754, 25261, 
    24606, 24030,
  27637, 27586, 27610, 27282, 26715, 25564, 24061, 23094, 22551, 22460, 
    22697, 23211, 24199, 25381, 26660, 27801, 27379, 26348, 25720, 25261, 
    24632, 24238,
  27560, 27540, 27462, 27188, 26601, 25550, 24064, 23099, 22592, 22469, 
    22740, 23180, 24132, 25293, 26095, 27619, 27149, 26269, 25734, 25310, 
    24670, 24151,
  27470, 27464, 27238, 27013, 26526, 25480, 24072, 23137, 22610, 22520, 
    22811, 23368, 24145, 25241, 26068, 27341, 26819, 25994, 25596, 25143, 
    24568, 24144,
  27373, 27363, 27101, 26867, 26412, 25443, 24057, 23111, 22603, 22514, 
    22779, 23386, 24155, 25290, 26385, 27091, 26351, 25828, 25444, 25118, 
    24529, 24063,
  27267, 27248, 26985, 26804, 26309, 25418, 24078, 23134, 22613, 22525, 
    22762, 23269, 24196, 25342, 26388, 26962, 26190, 25878, 25554, 25229, 
    24593, 24190,
  27151, 27119, 26919, 26681, 26282, 25365, 24002, 23119, 22580, 22588, 
    22785, 23284, 24063, 25297, 26517, 26882, 26401, 26051, 25713, 25229, 
    24631, 24103,
  27048, 26987, 26871, 26678, 26238, 25354, 24023, 23137, 22583, 22577, 
    22836, 23370, 24110, 25223, 26391, 26748, 26389, 26022, 25685, 25292, 
    24638, 24177,
  26988, 26895, 26815, 26640, 26240, 25357, 24040, 23128, 22574, 22557, 
    22756, 23291, 24265, 25460, 26662, 26712, 26246, 26051, 25685, 25204, 
    24612, 24251,
  26993, 26888, 26893, 26746, 26289, 25413, 24043, 23167, 22609, 22502, 
    22890, 23266, 24258, 25281, 26307, 26756, 26457, 26145, 25732, 25248, 
    24675, 24144,
  27052, 26958, 27025, 26813, 26332, 25379, 24102, 23146, 22670, 22548, 
    22796, 23286, 24184, 25286, 26644, 26840, 26607, 26189, 25823, 25285, 
    24663, 24177,
  27123, 27043, 27079, 26882, 26392, 25413, 24123, 23190, 22633, 22537, 
    22876, 23307, 24154, 25241, 26451, 26923, 26769, 26275, 25899, 25329, 
    24784, 24231,
  27159, 27091, 27054, 26932, 26400, 25483, 24130, 23137, 22641, 22591, 
    22833, 23360, 24334, 25318, 26100, 27032, 26912, 26304, 25892, 25360, 
    24784, 24337,
  27149, 27102, 27054, 26889, 26392, 25438, 24078, 23190, 22665, 22668, 
    22847, 23413, 24162, 25477, 26318, 26990, 26800, 26239, 25809, 25384, 
    24764, 24244,
  27128, 27110, 27003, 26851, 26360, 25348, 24064, 23234, 22633, 22594, 
    22765, 23294, 24206, 25346, 26531, 26809, 26526, 26124, 25726, 25254, 
    24771, 24231,
  27133, 27128, 26942, 26746, 26318, 25438, 24078, 23151, 22665, 22551, 
    22839, 23383, 24184, 25441, 26509, 26756, 26675, 26210, 25796, 25304, 
    24663, 24211,
  27159, 27138, 27023, 26832, 26385, 25438, 24082, 23184, 22680, 22674, 
    22853, 23309, 24120, 25337, 26307, 26821, 26650, 26260, 25775, 25267, 
    24631, 24056,
  27152, 27098, 27139, 26932, 26406, 25432, 24022, 23149, 22618, 22588, 
    22859, 23421, 24196, 25318, 26565, 26976, 26744, 26218, 25782, 25273, 
    24580, 24244,
  27042, 26962, 27154, 26982, 26429, 25410, 24067, 23193, 22650, 22632, 
    22842, 23357, 24241, 25246, 26157, 27093, 26663, 26232, 25768, 25198, 
    24638, 24063,
  26790, 26707, 27076, 26901, 26381, 25399, 24033, 23179, 22683, 22617, 
    22833, 23281, 24117, 25262, 26429, 27018, 26470, 26045, 25651, 25205, 
    24688, 24103,
  26441, 26377, 26810, 26703, 26320, 25368, 24099, 23196, 22677, 22660, 
    22944, 23335, 24212, 25313, 26187, 26748, 25997, 25647, 25526, 25062, 
    24561, 24084,
  26134, 26093, 26490, 26592, 26309, 25387, 24037, 23173, 22709, 22675, 
    22828, 23325, 24239, 25383, 26737, 26467, 25798, 25554, 25409, 25043, 
    24555, 24171,
  26031, 25995, 26528, 26535, 26246, 25365, 24050, 23155, 22735, 22612, 
    22785, 23363, 24229, 25248, 25882, 26426, 26339, 25835, 25485, 25068, 
    24536, 24077,
  26214, 26167, 26650, 26673, 26326, 25326, 24026, 23176, 22715, 22635, 
    22933, 23434, 24286, 25365, 26570, 26675, 26688, 26073, 25589, 25149, 
    24574, 24030,
  26622, 26587, 27076, 26945, 26460, 25405, 24006, 23170, 22701, 22635, 
    22802, 23376, 24056, 25288, 26291, 27224, 27235, 26319, 25726, 25242, 
    24645, 24111,
  27098, 27115, 27484, 27188, 26532, 25444, 24040, 23146, 22727, 22687, 
    22962, 23363, 24241, 25293, 26565, 27635, 27535, 26376, 25754, 25187, 
    24594, 24064,
  27484, 27566, 27569, 27235, 26572, 25410, 24020, 23191, 22684, 22690, 
    22939, 23315, 24180, 25407, 26197, 27812, 27635, 26493, 25838, 25193, 
    24594, 23990,
  27703, 27816, 27564, 27215, 26547, 25335, 23978, 23117, 22678, 22655, 
    22794, 23249, 24217, 25200, 26667, 27770, 27572, 26557, 25872, 25230, 
    24575, 24085,
  27776, 27867, 27498, 27188, 26554, 25382, 23999, 23144, 22713, 22707, 
    22863, 23280, 24276, 25253, 26479, 27706, 27660, 26601, 25948, 25243, 
    24575, 23951,
  27762, 27807, 27504, 27139, 26481, 25338, 23971, 23153, 22719, 22656, 
    22852, 23412, 24304, 25305, 26253, 27685, 27573, 26659, 25970, 25287, 
    24658, 24179,
  27704, 27720, 27485, 27172, 26487, 25360, 23912, 23144, 22716, 22713, 
    22943, 23402, 24161, 25335, 26557, 27647, 27510, 26651, 25990, 25318, 
    24550, 24159,
  27618, 27653, 27410, 27121, 26516, 25330, 23947, 23109, 22687, 22673, 
    22920, 23344, 24099, 25291, 26575, 27591, 27498, 26645, 25949, 25231, 
    24671, 24159,
  27521, 27610, 27326, 27075, 26401, 25274, 23906, 23104, 22676, 22737, 
    22921, 23501, 24361, 25338, 26485, 27497, 27529, 26681, 25997, 25287, 
    24595, 24099,
  27452, 27581, 27173, 27010, 26396, 25220, 23864, 23059, 22717, 22659, 
    22929, 23344, 24107, 25440, 26732, 27376, 27454, 26681, 26032, 25306, 
    24646, 24059,
  27442, 27558, 27115, 26929, 26250, 25193, 23805, 23057, 22694, 22700, 
    22918, 23464, 24208, 25447, 26573, 27265, 27310, 26667, 26079, 25318, 
    24621, 24119,
  27448, 27501, 27076, 26892, 26229, 25100, 23806, 23092, 22682, 22729, 
    22887, 23393, 24329, 25366, 26754, 27234, 27293, 26631, 25949, 25269, 
    24577, 23992,
  27291, 27268, 27072, 26798, 26164, 25117, 23837, 23057, 22685, 22764, 
    22916, 23388, 24391, 25420, 26735, 27226, 27094, 26371, 25853, 25182, 
    24462, 24087,
  26697, 26620, 27129, 26863, 26176, 25056, 23778, 23040, 22712, 22792, 
    22941, 23472, 24265, 25481, 26728, 27231, 27281, 26617, 26116, 25462, 
    24749, 24187,
  25490, 25399, 26948, 26731, 26124, 25058, 23778, 23069, 22709, 22790, 
    23016, 23409, 24241, 25574, 26343, 27175, 27448, 26826, 26219, 25524, 
    24743, 24114,
  23832, 23784, 25946, 26114, 25898, 24974, 23678, 23022, 22701, 22735, 
    22962, 23470, 24202, 25353, 26641, 26385, 27329, 26790, 26226, 25593, 
    24794, 24161,
  22292, 22353, 24088, 25064, 25452, 24846, 23674, 23034, 22771, 22745, 
    22962, 23389, 24345, 25509, 26724, 24193, 26148, 26682, 26295, 25704, 
    24909, 24309,
  21582, 21760, 22932, 24416, 25203, 24764, 23657, 23041, 22701, 22770, 
    23014, 23493, 24404, 25653, 26332, 22449, 25029, 26538, 26295, 25768, 
    25081, 24382,
  22072, 22276, 23614, 24798, 25298, 24768, 23650, 22976, 22716, 22791, 
    23074, 23547, 24304, 25604, 26750, 23095, 25247, 26610, 26337, 25867, 
    25113, 24497,
  23488, 23602, 25480, 25826, 25687, 24796, 23605, 23017, 22672, 22785, 
    23040, 23501, 24484, 25428, 26816, 25421, 26751, 26782, 26282, 25854, 
    25088, 24430,
  25104, 25109, 26684, 26504, 25876, 24815, 23582, 22950, 22755, 22768, 
    22946, 23469, 24366, 25514, 26564, 26918, 27356, 26820, 26365, 25793, 
    25063, 24544,
  26254, 26229, 26882, 26610, 25859, 24762, 23557, 23006, 22778, 22806, 
    22901, 23512, 24477, 25621, 26917, 27118, 27275, 26741, 26220, 25713, 
    25012, 24591,
  26685, 26704, 26854, 26562, 25801, 24692, 23513, 22935, 22734, 22780, 
    23027, 23644, 24339, 25714, 26876, 27085, 27281, 26662, 26131, 25526, 
    24942, 24484,
  26521, 26573, 26809, 26500, 25793, 24637, 23474, 22954, 22737, 22832, 
    22998, 23634, 24460, 25775, 26835, 27093, 27262, 26647, 26131, 25626, 
    24943, 24397,
  25994, 26022, 26745, 26449, 25719, 24637, 23475, 22972, 22729, 22824, 
    23081, 23568, 24507, 25663, 26749, 27009, 27225, 26632, 26145, 25552, 
    24937, 24351,
  25266, 25239, 26641, 26335, 25691, 24559, 23429, 22936, 22779, 22819, 
    23025, 23582, 24535, 25699, 26719, 26939, 27145, 26612, 26139, 25552, 
    24886, 24372,
  24422, 24380, 26264, 26172, 25542, 24533, 23402, 22913, 22782, 22827, 
    23028, 23516, 24444, 25726, 26809, 26601, 27170, 26612, 26167, 25559, 
    24829, 24365,
  23546, 23572, 25537, 25735, 25368, 24422, 23371, 22940, 22762, 22816, 
    23113, 23541, 24503, 25647, 27176, 25684, 26914, 26560, 26159, 25615, 
    24868, 24325,
  22745, 22885, 24888, 25367, 25256, 24369, 23330, 22955, 22786, 22894, 
    22963, 23623, 24565, 25645, 26854, 24461, 26268, 26489, 26063, 25578, 
    24874, 24319,
  22075, 22277, 24690, 25222, 25191, 24291, 23326, 22849, 22757, 22828, 
    23128, 23623, 24656, 25897, 27206, 23772, 26082, 26410, 26070, 25590, 
    24970, 24373,
  21449, 21608, 24701, 25266, 25093, 24243, 23271, 22861, 22760, 22871, 
    23034, 23565, 24674, 25764, 26698, 23554, 26132, 26432, 26091, 25659, 
    25008, 24400,
  20672, 20729, 24688, 25247, 25117, 24176, 23229, 22826, 22798, 22906, 
    23131, 23659, 24588, 25976, 26701, 23325, 26057, 26404, 26091, 25603, 
    25034, 24527,
  19704, 19666, 24630, 25220, 25051, 24151, 23185, 22841, 22755, 22904, 
    23243, 23644, 24707, 25825, 27157, 23207, 26157, 26389, 26016, 25486, 
    24945, 24487,
  18899, 18738, 24470, 25145, 24980, 24120, 23150, 22844, 22749, 22947, 
    23197, 23695, 24810, 25872, 26815, 23112, 26306, 26375, 25996, 25455, 
    24863, 24394,
  18728, 18328, 24526, 25148, 24960, 24081, 23091, 22783, 22820, 22861, 
    23146, 23764, 24618, 26154, 27139, 22933, 26485, 26238, 25803, 25343, 
    24615, 23940,
  19120, 18416, 24527, 25202, 24905, 23975, 23057, 22801, 22738, 22890, 
    23215, 23761, 24830, 26107, 26904, 22804, 26244, 26001, 25596, 24940, 
    24222, 23693,
  19393, 18543, 24747, 25197, 24886, 23841, 22998, 22769, 22794, 22950, 
    23280, 23855, 24828, 26270, 27159, 22676, 25269, 24949, 24708, 24351, 
    23790, 23345,
  28620, 28608, 27716, 26982, 25713, 24108, 22705, 22191, 22061, 22488, 
    22901, 23524, 24709, 25815, 26712, 28484, 28672, 27813, 27316, 26779, 
    25922, 25136,
  28581, 28571, 27759, 27109, 25850, 24242, 22735, 22223, 22069, 22445, 
    22878, 23625, 24509, 25660, 26314, 28548, 28765, 27856, 27351, 26748, 
    25954, 25089,
  28486, 28487, 27840, 27139, 25942, 24360, 22794, 22240, 22075, 22556, 
    22801, 23579, 24454, 25754, 26704, 28464, 28641, 27776, 27226, 26599, 
    25839, 25041,
  28381, 28405, 27663, 27150, 26025, 24477, 22895, 22287, 22080, 22384, 
    22812, 23422, 24439, 25801, 26422, 28288, 28498, 27690, 27171, 26679, 
    25807, 24954,
  28302, 28346, 27678, 27163, 26144, 24539, 22992, 22325, 22124, 22389, 
    22823, 23497, 24523, 25588, 26398, 28191, 28392, 27704, 27075, 26485, 
    25685, 24760,
  28271, 28315, 27657, 27214, 26144, 24648, 23040, 22337, 22124, 22449, 
    22715, 23449, 24397, 25623, 26548, 28201, 28335, 27697, 27101, 26468, 
    25628, 24807,
  28297, 28325, 27743, 27295, 26264, 24689, 23095, 22363, 22123, 22360, 
    22729, 23428, 24439, 25756, 26470, 28316, 28473, 27697, 27143, 26424, 
    25571, 24646,
  28368, 28383, 27929, 27413, 26370, 24821, 23178, 22439, 22146, 22475, 
    22851, 23393, 24345, 25704, 26248, 28484, 28691, 27726, 27067, 26399, 
    25469, 24378,
  28436, 28456, 27964, 27491, 26450, 24868, 23237, 22489, 22105, 22417, 
    22774, 23440, 24372, 25501, 26179, 28601, 28709, 27718, 26991, 26225, 
    25322, 24465,
  28450, 28491, 28065, 27569, 26504, 24941, 23271, 22477, 22163, 22397, 
    22725, 23440, 24270, 25650, 26407, 28548, 28647, 27581, 26853, 26088, 
    25131, 24244,
  28403, 28463, 27931, 27482, 26526, 24949, 23323, 22464, 22168, 22356, 
    22787, 23366, 24334, 25503, 26503, 28470, 28566, 27523, 26667, 25914, 
    24914, 23996,
  28324, 28388, 27847, 27401, 26490, 25022, 23365, 22509, 22162, 22427, 
    22750, 23394, 24299, 25624, 26485, 28285, 28348, 27379, 26598, 25771, 
    24761, 23975,
  28238, 28282, 27763, 27367, 26532, 25061, 23379, 22585, 22168, 22378, 
    22704, 23343, 24200, 25436, 26370, 28182, 28335, 27472, 26729, 25770, 
    24818, 24089,
  28139, 28156, 27771, 27394, 26596, 25145, 23493, 22611, 22220, 22421, 
    22750, 23310, 24279, 25379, 26365, 28194, 28460, 27624, 26845, 25957, 
    24869, 24122,
  28024, 28027, 27784, 27364, 26567, 25201, 23496, 22640, 22176, 22470, 
    22775, 23310, 24195, 25384, 26585, 28096, 28367, 27588, 26790, 25869, 
    24913, 24135,
  27920, 27934, 27626, 27324, 26598, 25204, 23562, 22672, 22217, 22423, 
    22749, 23444, 24252, 25338, 26932, 27907, 28110, 27429, 26651, 25832, 
    24957, 24155,
  27868, 27901, 27429, 27197, 26501, 25156, 23565, 22654, 22205, 22406, 
    22709, 23342, 24217, 25377, 26674, 27740, 27894, 27184, 26438, 25676, 
    24855, 24188,
  27878, 27918, 27515, 27232, 26592, 25273, 23666, 22734, 22260, 22377, 
    22777, 23378, 24224, 25281, 26345, 27782, 27906, 27132, 26279, 25521, 
    24817, 24214,
  27926, 27958, 27674, 27437, 26654, 25365, 23686, 22752, 22286, 22414, 
    22779, 23332, 24327, 25521, 26604, 28032, 28037, 26981, 26238, 25552, 
    24867, 24227,
  27973, 28007, 27810, 27463, 26747, 25382, 23728, 22825, 22286, 22382, 
    22774, 23435, 24283, 25318, 26309, 28154, 28049, 26794, 26024, 25421, 
    24772, 24214,
  27994, 28049, 27824, 27466, 26760, 25419, 23772, 22822, 22315, 22413, 
    22890, 23336, 24189, 25453, 26548, 28172, 27999, 26692, 25989, 25309, 
    24606, 24100,
  27995, 28073, 27796, 27485, 26698, 25432, 23758, 22827, 22323, 22410, 
    22773, 23219, 24137, 25590, 26118, 28097, 27900, 26626, 25954, 25346, 
    24669, 23985,
  27986, 28060, 27682, 27347, 26672, 25390, 23810, 22865, 22358, 22399, 
    22721, 23343, 24174, 25486, 26420, 27979, 27701, 26626, 25947, 25364, 
    24650, 24065,
  27940, 27970, 27585, 27279, 26629, 25399, 23821, 22874, 22341, 22464, 
    22747, 23366, 24173, 25231, 26790, 27868, 27495, 26497, 25906, 25358, 
    24681, 24152,
  27799, 27746, 27575, 27342, 26615, 25396, 23855, 22912, 22346, 22401, 
    22781, 23325, 24099, 25264, 26369, 27907, 27520, 26497, 25857, 25351, 
    24656, 24018,
  27535, 27386, 27582, 27326, 26682, 25454, 23858, 22915, 22387, 22389, 
    22707, 23287, 24148, 25329, 26231, 27894, 27564, 26468, 25891, 25289, 
    24636, 24045,
  27203, 26986, 27301, 27151, 26589, 25407, 23851, 22947, 22422, 22435, 
    22695, 23383, 24074, 25201, 26216, 27651, 27526, 26439, 25843, 25295, 
    24687, 24071,
  26925, 26693, 26979, 26962, 26534, 25437, 23886, 22923, 22454, 22415, 
    22815, 23299, 24116, 25420, 26407, 27317, 27307, 26396, 25822, 25282, 
    24680, 24044,
  26809, 26592, 26870, 26929, 26479, 25418, 23942, 22970, 22430, 22423, 
    22740, 23339, 24192, 25196, 26579, 27189, 27226, 26323, 25807, 25288, 
    24642, 24064,
  26877, 26676, 27020, 27010, 26543, 25490, 23959, 22970, 22433, 22400, 
    22754, 23306, 24076, 25163, 26545, 27335, 27282, 26272, 25746, 25207, 
    24610, 23990,
  27048, 26866, 27225, 27126, 26597, 25524, 24021, 23041, 22485, 22451, 
    22674, 23240, 24266, 25072, 26221, 27534, 27296, 26316, 25779, 25151, 
    24622, 24030,
  27211, 27065, 27304, 27137, 26614, 25476, 23962, 22990, 22479, 22459, 
    22668, 23364, 24191, 25056, 26247, 27537, 27264, 26287, 25738, 25163, 
    24609, 24097,
  27307, 27192, 27164, 27073, 26620, 25512, 23972, 23029, 22473, 22445, 
    22793, 23390, 24120, 25289, 26460, 27432, 27126, 26207, 25690, 25126, 
    24552, 23976,
  27345, 27230, 27162, 27094, 26582, 25493, 24031, 23029, 22491, 22453, 
    22745, 23321, 24110, 25242, 26499, 27443, 27096, 26149, 25654, 25194, 
    24596, 24003,
  27354, 27222, 27248, 27134, 26631, 25532, 23993, 23034, 22520, 22445, 
    22751, 23351, 24122, 25328, 26400, 27549, 26996, 26076, 25635, 25150, 
    24532, 24103,
  27343, 27212, 27319, 27179, 26625, 25495, 24024, 23117, 22508, 22444, 
    22716, 23313, 24043, 25196, 26097, 27624, 26947, 26054, 25586, 25088, 
    24468, 24062,
  27306, 27203, 27299, 27150, 26539, 25501, 24031, 23134, 22543, 22444, 
    22787, 23252, 24193, 25249, 26421, 27563, 26754, 26012, 25593, 25076, 
    24519, 24062,
  27245, 27173, 27220, 27016, 26534, 25495, 24038, 23116, 22522, 22533, 
    22705, 23244, 24048, 25191, 26710, 27343, 26585, 26026, 25586, 25156, 
    24538, 24022,
  27165, 27105, 27106, 26918, 26425, 25420, 24055, 23060, 22540, 22430, 
    22730, 23259, 24114, 25440, 26356, 27048, 26349, 25881, 25558, 25138, 
    24564, 23968,
  27066, 27001, 26923, 26695, 26304, 25374, 23989, 23086, 22569, 22435, 
    22710, 23231, 24035, 25253, 26416, 26704, 25863, 25672, 25434, 25156, 
    24538, 24049,
  26938, 26870, 26814, 26573, 26235, 25321, 24010, 23137, 22519, 22444, 
    22730, 23208, 24141, 25142, 26035, 26529, 25632, 25665, 25496, 25050, 
    24480, 23955,
  26791, 26723, 26712, 26598, 26126, 25304, 24030, 23113, 22601, 22449, 
    22775, 23294, 24107, 25223, 26095, 26460, 25938, 25851, 25606, 25168, 
    24653, 23995,
  26660, 26585, 26603, 26528, 26141, 25318, 24017, 23113, 22595, 22550, 
    22787, 23269, 24102, 24985, 26240, 26416, 26062, 25881, 25626, 25069, 
    24500, 24095,
  26590, 26507, 26641, 26515, 26247, 25304, 24034, 23131, 22598, 22536, 
    22787, 23221, 24013, 25260, 26335, 26401, 25664, 25787, 25565, 25168, 
    24620, 24082,
  26608, 26529, 26710, 26593, 26245, 25304, 24065, 23157, 22569, 22504, 
    22715, 23256, 24141, 25253, 26525, 26424, 25788, 25794, 25599, 25093, 
    24570, 24061,
  26705, 26634, 26801, 26684, 26256, 25374, 24037, 23145, 22589, 22492, 
    22827, 23274, 24205, 25227, 26360, 26560, 26038, 25874, 25620, 25224, 
    24640, 24082,
  26833, 26758, 26943, 26785, 26329, 25430, 24037, 23139, 22610, 22484, 
    22704, 23350, 24064, 25340, 26201, 26710, 25938, 25801, 25530, 25193, 
    24595, 24028,
  26932, 26850, 26968, 26826, 26326, 25400, 24051, 23125, 22607, 22510, 
    22801, 23269, 24205, 25372, 26244, 26725, 25925, 25831, 25551, 25187, 
    24627, 24108,
  26979, 26902, 26951, 26797, 26335, 25358, 24037, 23193, 22648, 22461, 
    22727, 23251, 23988, 25330, 26429, 26707, 26168, 26018, 25682, 25255, 
    24729, 24142,
  26989, 26929, 26882, 26746, 26316, 25360, 24016, 23178, 22598, 22467, 
    22707, 23251, 24180, 25181, 26341, 26601, 26118, 25917, 25675, 25187, 
    24608, 24156,
  26982, 26934, 26826, 26743, 26287, 25352, 24030, 23181, 22636, 22550, 
    22815, 23310, 24027, 25337, 26507, 26457, 25714, 25607, 25454, 25156, 
    24665, 24122,
  26950, 26902, 26938, 26749, 26342, 25405, 24044, 23163, 22616, 22561, 
    22767, 23282, 24245, 25321, 26324, 26557, 25645, 25685, 25461, 25112, 
    24633, 24109,
  26857, 26806, 26994, 26826, 26332, 25397, 24058, 23139, 22645, 22619, 
    22804, 23287, 24030, 25099, 26576, 26803, 26087, 25729, 25496, 25119, 
    24576, 24089,
  26660, 26608, 26904, 26810, 26347, 25352, 24023, 23157, 22653, 22570, 
    22861, 23244, 24109, 25358, 26528, 26881, 26044, 25650, 25440, 25094, 
    24474, 23968,
  26340, 26287, 26771, 26651, 26301, 25338, 23992, 23184, 22645, 22547, 
    22832, 23251, 24233, 25316, 26379, 26654, 25857, 25607, 25385, 25087, 
    24480, 24015,
  25950, 25897, 26464, 26474, 26242, 25290, 24020, 23140, 22680, 22547, 
    22850, 23269, 24112, 25318, 26491, 26340, 25484, 25441, 25302, 25025, 
    24519, 23961,
  25628, 25578, 26238, 26329, 26176, 25344, 24010, 23146, 22619, 22584, 
    22824, 23315, 24124, 25244, 26282, 26123, 25969, 25737, 25496, 25131, 
    24564, 24109,
  25541, 25499, 26060, 26296, 26150, 25279, 23999, 23110, 22607, 22585, 
    22881, 23279, 24265, 25221, 26132, 26087, 26329, 25954, 25572, 25125, 
    24653, 23975,
  25782, 25749, 26324, 26428, 26182, 25333, 23940, 23160, 22642, 22617, 
    22816, 23275, 24159, 25351, 26537, 26374, 26822, 26235, 25710, 25281, 
    24697, 24136,
  26293, 26278, 26826, 26798, 26416, 25397, 23965, 23137, 22689, 22662, 
    22776, 23399, 24285, 25153, 26431, 26978, 27239, 26451, 25882, 25324, 
    24583, 24096,
  26895, 26918, 27316, 27042, 26491, 25375, 23944, 23137, 22663, 22651, 
    22856, 23333, 24048, 25498, 26329, 27554, 27569, 26518, 25869, 25250, 
    24609, 24116,
  27394, 27469, 27547, 27237, 26562, 25406, 23965, 23143, 22684, 22617, 
    22804, 23295, 24122, 25419, 26388, 27772, 27650, 26604, 25890, 25250, 
    24545, 24130,
  27686, 27801, 27560, 27229, 26537, 25339, 23944, 23143, 22684, 22634, 
    22885, 23260, 24347, 25403, 26071, 27763, 27582, 26632, 25918, 25306, 
    24565, 24049,
  27785, 27908, 27484, 27191, 26525, 25344, 23934, 23117, 22684, 22623, 
    22885, 23313, 24295, 25349, 26457, 27721, 27669, 26698, 26063, 25306, 
    24590, 24090,
  27774, 27877, 27453, 27169, 26485, 25339, 23938, 23100, 22708, 22669, 
    22916, 23395, 24308, 25387, 26468, 27699, 27582, 26698, 26035, 25288, 
    24667, 24090,
  27723, 27809, 27501, 27081, 26471, 25302, 23886, 23091, 22676, 22718, 
    22840, 23362, 24103, 25303, 26421, 27707, 27675, 26785, 26056, 25325, 
    24635, 24110,
  27658, 27754, 27501, 27148, 26422, 25322, 23882, 23100, 22696, 22655, 
    22879, 23454, 24263, 25443, 26492, 27671, 27769, 26785, 26070, 25369, 
    24635, 24071,
  27581, 27712, 27404, 27118, 26434, 25302, 23872, 23082, 22688, 22715, 
    22808, 23347, 24145, 25322, 26146, 27587, 27756, 26843, 26098, 25431, 
    24661, 24145,
  27499, 27655, 27299, 26989, 26357, 25210, 23869, 23079, 22673, 22684, 
    22811, 23261, 24301, 25553, 26700, 27417, 27532, 26885, 26195, 25419, 
    24655, 24158,
  27426, 27556, 27164, 26922, 26288, 25185, 23844, 23080, 22685, 22661, 
    23008, 23352, 24282, 25250, 26685, 27328, 27414, 26865, 26222, 25463, 
    24738, 24192,
  27312, 27366, 27063, 26844, 26245, 25109, 23803, 23033, 22706, 22693, 
    22969, 23368, 24207, 25341, 26603, 27257, 27326, 26771, 26174, 25351, 
    24655, 24005,
  26978, 26954, 27053, 26809, 26156, 25062, 23754, 23048, 22691, 22691, 
    22920, 23302, 24245, 25353, 26466, 27174, 27301, 26750, 26209, 25507, 
    24770, 24172,
  26162, 26109, 26959, 26739, 26145, 25051, 23779, 23077, 22700, 22682, 
    22849, 23386, 24368, 25369, 26749, 27196, 27371, 26829, 26244, 25637, 
    24745, 24159,
  24725, 24704, 26409, 26437, 25948, 25015, 23741, 23037, 22709, 22700, 
    22967, 23404, 24321, 25810, 26616, 26873, 27401, 26857, 26306, 25694, 
    24873, 24226,
  22891, 22950, 25040, 25555, 25650, 24902, 23675, 23031, 22678, 22746, 
    22907, 23506, 24240, 25423, 26410, 25452, 26985, 26894, 26341, 25688, 
    24956, 24240,
  21296, 21457, 23225, 24583, 25259, 24765, 23651, 22998, 22716, 22740, 
    22981, 23460, 24196, 25567, 26604, 23153, 25517, 26657, 26320, 25806, 
    25026, 24367,
  20678, 20901, 22397, 24139, 25104, 24754, 23647, 22990, 22701, 22683, 
    22905, 23491, 24413, 25491, 26710, 21713, 24920, 26606, 26299, 25837, 
    25115, 24368,
  21368, 21542, 23383, 24683, 25316, 24738, 23634, 22999, 22725, 22747, 
    22919, 23509, 24275, 25549, 26632, 22618, 25225, 26678, 26314, 25738, 
    25109, 24435,
  22994, 23025, 25453, 25778, 25645, 24797, 23600, 22979, 22801, 22741, 
    22993, 23469, 24401, 25440, 26756, 25270, 26817, 26785, 26307, 25732, 
    25116, 24602,
  24724, 24632, 26663, 26500, 25876, 24791, 23600, 22976, 22752, 22753, 
    23013, 23532, 24293, 25586, 26645, 26928, 27396, 26787, 26328, 25850, 
    25224, 24616,
  25832, 25731, 26891, 26567, 25866, 24763, 23565, 22988, 22796, 22776, 
    23002, 23462, 24587, 25675, 26648, 27134, 27265, 26751, 26266, 25726, 
    25097, 24590,
  26090, 26059, 26787, 26507, 25746, 24671, 23496, 22956, 22755, 22808, 
    22977, 23480, 24456, 25484, 26476, 27076, 27235, 26765, 26266, 25789, 
    25161, 24623,
  25700, 25724, 26635, 26419, 25720, 24590, 23500, 22986, 22747, 22799, 
    23071, 23460, 24397, 25676, 26597, 26994, 27154, 26723, 26225, 25707, 
    25060, 24584,
  24983, 25002, 26506, 26309, 25646, 24565, 23458, 22924, 22756, 22811, 
    23012, 23523, 24356, 25692, 26588, 26857, 27135, 26665, 26218, 25721, 
    24964, 24537,
  24158, 24151, 26304, 26116, 25600, 24484, 23445, 22924, 22753, 22849, 
    23020, 23521, 24573, 25690, 26528, 26648, 27110, 26571, 26184, 25659, 
    24965, 24263,
  23339, 23347, 25607, 25793, 25437, 24456, 23358, 22936, 22780, 22832, 
    22984, 23600, 24556, 25813, 26657, 25935, 26910, 26564, 26122, 25678, 
    24965, 24364,
  22619, 22707, 24720, 25360, 25272, 24389, 23362, 22925, 22768, 22824, 
    22970, 23608, 24653, 25651, 26487, 24562, 26332, 26521, 26087, 25591, 
    24965, 24324,
  22092, 22269, 24510, 25115, 25201, 24336, 23307, 22910, 22780, 22841, 
    23050, 23575, 24589, 25857, 26704, 23605, 25810, 26499, 26109, 25635, 
    24972, 24458,
  21757, 21949, 24710, 25252, 25172, 24250, 23328, 22866, 22775, 22816, 
    23047, 23598, 24539, 25816, 26741, 23607, 26072, 26493, 26135, 25772, 
    24947, 24425,
  21440, 21552, 24799, 25314, 25118, 24241, 23286, 22852, 22784, 22839, 
    23042, 23659, 24461, 25851, 26956, 23637, 26060, 26535, 26157, 25846, 
    25119, 24639,
  20878, 20881, 24797, 25290, 25118, 24163, 23227, 22841, 22775, 22870, 
    23150, 23614, 24653, 26029, 27129, 23483, 26110, 26471, 26109, 25648, 
    25094, 24552,
  19997, 19935, 24743, 25269, 25035, 24138, 23176, 22835, 22723, 22851, 
    23114, 23675, 24676, 25865, 26753, 23365, 26247, 26464, 26060, 25530, 
    25011, 24600,
  19142, 19003, 24470, 25177, 24984, 24043, 23117, 22850, 22750, 22842, 
    23026, 23736, 24656, 25926, 26548, 23016, 26297, 26435, 26060, 25604, 
    24942, 24440,
  18809, 18458, 24455, 25130, 24961, 24013, 23100, 22797, 22796, 22829, 
    23159, 23671, 24644, 26121, 26942, 22592, 26328, 26328, 25957, 25382, 
    24720, 24199,
  19011, 18355, 24562, 25105, 24873, 23904, 23031, 22809, 22753, 22889, 
    23157, 23818, 24738, 26038, 26982, 22368, 26160, 26176, 25724, 25128, 
    24421, 23778,
  19197, 18389, 24676, 25146, 24879, 23837, 23013, 22765, 22747, 22895, 
    23203, 23714, 24893, 25989, 26645, 22295, 25651, 25463, 25070, 24606, 
    24052, 23525,
  28624, 28639, 27751, 27044, 25753, 24128, 22703, 22193, 22097, 22470, 
    22905, 23625, 24476, 25799, 26672, 28485, 28687, 27869, 27322, 26754, 
    25929, 25099,
  28583, 28603, 27803, 27132, 25828, 24229, 22755, 22187, 22062, 22455, 
    22807, 23554, 24609, 25689, 26691, 28495, 28724, 27775, 27294, 26742, 
    25873, 24999,
  28485, 28520, 27835, 27154, 25982, 24343, 22838, 22239, 22085, 22418, 
    22801, 23498, 24444, 25838, 26257, 28495, 28662, 27782, 27197, 26654, 
    25751, 24852,
  28380, 28435, 27759, 27165, 26035, 24461, 22938, 22271, 22102, 22446, 
    22787, 23554, 24481, 25729, 26800, 28329, 28475, 27659, 27107, 26537, 
    25713, 24838,
  28302, 28368, 27722, 27126, 26081, 24550, 22948, 22315, 22082, 22454, 
    22738, 23543, 24296, 25530, 26899, 28216, 28432, 27667, 27079, 26474, 
    25649, 24797,
  28264, 28323, 27682, 27181, 26160, 24635, 23055, 22365, 22117, 22417, 
    22732, 23538, 24330, 25717, 26250, 28160, 28313, 27753, 27079, 26499, 
    25649, 24737,
  28278, 28315, 27785, 27278, 26282, 24702, 23125, 22365, 22134, 22419, 
    22863, 23462, 24493, 25610, 26528, 28224, 28450, 27746, 27114, 26424, 
    25534, 24717,
  28336, 28359, 27950, 27379, 26332, 24805, 23183, 22423, 22183, 22410, 
    22817, 23451, 24260, 25547, 26521, 28366, 28599, 27760, 27059, 26354, 
    25483, 24555,
  28400, 28431, 27960, 27429, 26426, 24911, 23246, 22485, 22145, 22441, 
    22709, 23469, 24408, 25507, 26613, 28464, 28581, 27645, 26921, 26244, 
    25298, 24462,
  28415, 28473, 27970, 27507, 26490, 24987, 23283, 22494, 22165, 22476, 
    22780, 23395, 24400, 25427, 26724, 28476, 28649, 27579, 26851, 26038, 
    25063, 24100,
  28361, 28446, 27881, 27488, 26553, 25017, 23384, 22567, 22162, 22415, 
    22771, 23438, 24299, 25416, 26559, 28342, 28487, 27500, 26782, 25895, 
    24973, 24066,
  28267, 28362, 27876, 27429, 26559, 25014, 23415, 22558, 22191, 22438, 
    22771, 23417, 24343, 25629, 26390, 28235, 28518, 27579, 26810, 26050, 
    24992, 24059,
  28168, 28252, 27785, 27472, 26564, 25070, 23484, 22628, 22214, 22412, 
    22784, 23478, 24314, 25474, 26554, 28197, 28407, 27629, 26941, 26087, 
    25074, 24273,
  28073, 28130, 27762, 27409, 26570, 25162, 23498, 22622, 22245, 22417, 
    22762, 23371, 24348, 25408, 26910, 28179, 28456, 27644, 27003, 26179, 
    25157, 24306,
  27979, 28010, 27704, 27375, 26526, 25202, 23504, 22684, 22181, 22405, 
    22747, 23348, 24222, 25352, 26566, 28051, 28282, 27500, 26775, 25938, 
    25010, 24279,
  27900, 27924, 27574, 27297, 26554, 25204, 23580, 22710, 22251, 22411, 
    22735, 23348, 24199, 25334, 26885, 27867, 28057, 27196, 26401, 25657, 
    24870, 24232,
  27867, 27898, 27546, 27256, 26535, 25251, 23577, 22751, 22324, 22416, 
    22823, 23304, 24263, 25424, 26595, 27735, 27871, 27001, 26244, 25564, 
    24888, 24419,
  27893, 27923, 27572, 27276, 26578, 25302, 23674, 22733, 22265, 22470, 
    22749, 23444, 24191, 25393, 26549, 27803, 27826, 26835, 26174, 25546, 
    24844, 24285,
  27951, 27965, 27759, 27442, 26690, 25347, 23667, 22774, 22268, 22444, 
    22746, 23395, 24098, 25142, 26151, 28088, 28045, 26821, 26160, 25458, 
    24844, 24204,
  27997, 28000, 27914, 27571, 26778, 25394, 23767, 22830, 22317, 22478, 
    22749, 23352, 24302, 25424, 26482, 28207, 28057, 26647, 25953, 25427, 
    24766, 24211,
  28003, 28016, 27826, 27482, 26754, 25369, 23757, 22835, 22308, 22490, 
    22703, 23371, 24205, 25372, 26546, 28119, 27907, 26604, 25967, 25290, 
    24728, 24183,
  27975, 28007, 27651, 27379, 26657, 25363, 23781, 22829, 22392, 22446, 
    22725, 23377, 24230, 25542, 26495, 27932, 27578, 26460, 25863, 25320, 
    24671, 24090,
  27925, 27960, 27589, 27272, 26626, 25352, 23812, 22891, 22354, 22423, 
    22756, 23313, 24289, 25293, 26635, 27762, 27404, 26379, 25828, 25289, 
    24651, 24096,
  27841, 27844, 27548, 27269, 26603, 25366, 23808, 22897, 22383, 22434, 
    22790, 23280, 24215, 25263, 26401, 27715, 27323, 26387, 25835, 25301, 
    24651, 24096,
  27683, 27615, 27589, 27328, 26637, 25410, 23867, 22946, 22392, 22480, 
    22710, 23318, 24131, 25437, 26524, 27787, 27316, 26423, 25869, 25307, 
    24689, 24028,
  27443, 27280, 27451, 27291, 26675, 25469, 23846, 22914, 22430, 22451, 
    22824, 23322, 24177, 25484, 26160, 27748, 27379, 26357, 25793, 25251, 
    24625, 24048,
  27168, 26934, 27142, 27101, 26632, 25438, 23877, 22987, 22406, 22439, 
    22744, 23396, 24175, 25169, 26351, 27447, 27173, 26271, 25731, 25232, 
    24631, 24048,
  26946, 26700, 26800, 26894, 26517, 25435, 23915, 22990, 22441, 22479, 
    22846, 23309, 24160, 25360, 26594, 27141, 27148, 26285, 25731, 25232, 
    24612, 24001,
  26849, 26637, 26850, 26951, 26543, 25477, 23915, 23013, 22447, 22447, 
    22749, 23284, 24103, 25132, 26417, 27082, 26992, 26104, 25710, 25182, 
    24573, 24047,
  26883, 26706, 27109, 27060, 26582, 25519, 23950, 23010, 22423, 22502, 
    22772, 23235, 24172, 25260, 26390, 27266, 26812, 26032, 25530, 25170, 
    24547, 23913,
  26981, 26821, 27299, 27135, 26610, 25533, 23939, 23016, 22502, 22476, 
    22774, 23342, 24134, 25276, 26307, 27375, 26625, 25823, 25468, 25082, 
    24516, 24107,
  27058, 26906, 27287, 27128, 26617, 25496, 23953, 23028, 22476, 22516, 
    22774, 23291, 24162, 25227, 26184, 27325, 26457, 25765, 25406, 25001, 
    24477, 23986,
  27077, 26923, 27129, 27026, 26591, 25485, 24016, 23063, 22540, 22478, 
    22763, 23412, 24157, 25429, 26494, 27178, 26351, 25657, 25364, 25007, 
    24509, 23933,
  27059, 26890, 27015, 26975, 26534, 25468, 23998, 23096, 22557, 22418, 
    22771, 23331, 24062, 25226, 26112, 27119, 26345, 25714, 25378, 24970, 
    24420, 23799,
  27032, 26854, 27013, 26975, 26520, 25499, 24005, 23110, 22540, 22498, 
    22739, 23295, 24211, 25247, 26274, 27122, 26388, 25785, 25488, 25076, 
    24521, 23986,
  27007, 26843, 26923, 26859, 26514, 25507, 24012, 23119, 22539, 22523, 
    22757, 23287, 24280, 25170, 26266, 27054, 26438, 25945, 25550, 25132, 
    24534, 23959,
  26973, 26841, 26997, 26862, 26468, 25437, 24025, 23104, 22557, 22512, 
    22745, 23280, 24082, 25380, 26622, 27007, 26407, 25945, 25578, 25156, 
    24559, 24106,
  26920, 26816, 26939, 26862, 26413, 25443, 24036, 23101, 22562, 22520, 
    22776, 23249, 24099, 25438, 26300, 26960, 26463, 26068, 25660, 25156, 
    24591, 23985,
  26838, 26742, 26954, 26789, 26376, 25404, 24018, 23124, 22580, 22478, 
    22759, 23267, 24126, 25252, 26387, 26791, 26276, 26003, 25604, 25087, 
    24521, 24066,
  26709, 26609, 26870, 26710, 26301, 25364, 24042, 23145, 22580, 22586, 
    22748, 23353, 24163, 25270, 26457, 26482, 25728, 25857, 25536, 25143, 
    24539, 24153,
  26530, 26429, 26698, 26538, 26204, 25358, 24018, 23121, 22597, 22469, 
    22819, 23262, 24022, 25198, 26207, 26301, 25603, 25707, 25474, 25081, 
    24571, 24146,
  26325, 26232, 26532, 26449, 26129, 25288, 24066, 23165, 22588, 22457, 
    22782, 23203, 24217, 25469, 26247, 26279, 25734, 25793, 25584, 25143, 
    24609, 24132,
  26152, 26067, 26487, 26425, 26167, 25364, 24028, 23186, 22635, 22508, 
    22813, 23284, 24190, 25270, 26353, 26243, 25826, 25865, 25543, 25075, 
    24629, 24058,
  26066, 25985, 26388, 26403, 26179, 25383, 24049, 23177, 22644, 22609, 
    22753, 23254, 24165, 25450, 26167, 26145, 25578, 25670, 25480, 25162, 
    24603, 24079,
  26091, 26015, 26396, 26422, 26164, 25372, 24053, 23156, 22626, 22503, 
    22727, 23416, 24187, 25098, 26260, 26117, 25329, 25641, 25459, 25149, 
    24654, 24079,
  26212, 26135, 26589, 26557, 26242, 25369, 24042, 23147, 22632, 22554, 
    22770, 23259, 24178, 25214, 26312, 26268, 25815, 25713, 25563, 25162, 
    24629, 24092,
  26377, 26290, 26731, 26646, 26299, 25420, 24074, 23183, 22632, 22549, 
    22824, 23294, 24039, 25247, 26151, 26321, 25771, 25678, 25522, 25187, 
    24603, 24099,
  26528, 26430, 26785, 26743, 26273, 25412, 24042, 23212, 22652, 22574, 
    22858, 23320, 24316, 25268, 26260, 26396, 25715, 25735, 25556, 25149, 
    24609, 24139,
  26633, 26529, 26819, 26724, 26287, 25372, 24091, 23186, 22632, 22600, 
    22812, 23368, 24042, 25317, 26295, 26443, 25771, 25750, 25528, 25218, 
    24629, 24199,
  26687, 26580, 26804, 26694, 26307, 25403, 24035, 23203, 22638, 22571, 
    22853, 23305, 24128, 25163, 26454, 26401, 25435, 25446, 25273, 25037, 
    24565, 24058,
  26681, 26577, 26817, 26756, 26293, 25392, 24025, 23171, 22685, 22569, 
    22864, 23335, 24225, 25329, 26072, 26399, 24794, 24926, 25011, 24863, 
    24469, 24099,
  26599, 26515, 26832, 26692, 26256, 25414, 24039, 23168, 22682, 22606, 
    22844, 23343, 23992, 25121, 26373, 26415, 24794, 24984, 25059, 24944, 
    24450, 23945,
  26426, 26377, 26746, 26700, 26287, 25395, 24025, 23198, 22647, 22589, 
    22787, 23315, 24126, 25296, 26520, 26499, 25086, 25100, 25135, 24913, 
    24545, 24065,
  26156, 26133, 26581, 26598, 26247, 25398, 24022, 23209, 22655, 22563, 
    22873, 23267, 24165, 25149, 26254, 26407, 25186, 25093, 25122, 24906, 
    24450, 24045,
  25795, 25772, 26388, 26476, 26224, 25344, 24049, 23183, 22723, 22626, 
    22804, 23267, 24163, 25314, 26378, 26215, 25124, 25013, 24983, 24826, 
    24361, 23905,
  25393, 25350, 26134, 26366, 26196, 25291, 24001, 23142, 22650, 22638, 
    22850, 23391, 24054, 25340, 26390, 25992, 25417, 25244, 25149, 24926, 
    24475, 24086,
  25074, 25014, 25929, 26225, 26165, 25291, 24046, 23169, 22706, 22666, 
    22916, 23445, 24035, 25513, 26240, 25757, 26082, 25764, 25446, 25112, 
    24476, 24119,
  25001, 24947, 25776, 26139, 26104, 25347, 24011, 23180, 22691, 22678, 
    22944, 23351, 24089, 25391, 26557, 25626, 26469, 26068, 25598, 25150, 
    24540, 24006,
  25279, 25249, 26004, 26242, 26135, 25373, 24012, 23148, 22662, 22635, 
    22807, 23414, 24220, 25312, 26470, 25897, 26743, 26349, 25840, 25274, 
    24706, 24126,
  25869, 25867, 26497, 26598, 26293, 25350, 23966, 23151, 22671, 22658, 
    22999, 23409, 24193, 25301, 26475, 26526, 27142, 26516, 25867, 25268, 
    24648, 24139,
  26592, 26619, 27175, 26982, 26468, 25387, 23984, 23181, 22718, 22604, 
    22813, 23318, 24166, 25268, 26285, 27301, 27490, 26566, 25923, 25287, 
    24636, 24073,
  27227, 27292, 27520, 27188, 26531, 25378, 23949, 23157, 22650, 22647, 
    22908, 23321, 24196, 25254, 26603, 27665, 27671, 26631, 25937, 25281, 
    24655, 24093,
  27631, 27743, 27535, 27174, 26510, 25342, 23925, 23089, 22659, 22670, 
    22871, 23415, 24159, 25371, 26453, 27721, 27640, 26754, 26034, 25380, 
    24706, 24154,
  27795, 27944, 27441, 27179, 26500, 25334, 23970, 23143, 22706, 22579, 
    22823, 23392, 24218, 25406, 26499, 27660, 27671, 26790, 26103, 25406, 
    24732, 24100,
  27807, 27968, 27454, 27156, 26471, 25348, 23925, 23125, 22678, 22665, 
    22920, 23364, 24041, 25525, 26610, 27604, 27651, 26906, 26096, 25481, 
    24681, 24187,
  27765, 27914, 27421, 27172, 26457, 25303, 23943, 23164, 22684, 22634, 
    22803, 23385, 24169, 25597, 26431, 27640, 27696, 26899, 26151, 25568, 
    24675, 24208,
  27704, 27833, 27393, 27123, 26434, 25345, 23894, 23114, 22704, 22703, 
    22854, 23319, 24312, 25343, 26473, 27576, 27676, 26863, 26193, 25580, 
    24821, 24208,
  27602, 27719, 27332, 27091, 26394, 25270, 23891, 23114, 22669, 22697, 
    22963, 23339, 24236, 25446, 26342, 27584, 27721, 26921, 26248, 25606, 
    24866, 24262,
  27431, 27538, 27241, 26964, 26357, 25247, 23888, 23102, 22754, 22734, 
    22909, 23520, 24273, 25383, 26417, 27484, 27640, 26935, 26166, 25512, 
    24797, 24235,
  27191, 27272, 27163, 26954, 26301, 25174, 23849, 23100, 22728, 22729, 
    22918, 23401, 24237, 25372, 26785, 27353, 27491, 26820, 26173, 25500, 
    24790, 24202,
  26858, 26899, 27092, 26857, 26260, 25183, 23812, 23067, 22740, 22732, 
    22921, 23426, 24335, 25444, 26629, 27289, 27441, 26842, 26145, 25681, 
    24835, 24269,
  26313, 26332, 27035, 26776, 26159, 25034, 23753, 23056, 22775, 22729, 
    22972, 23399, 24168, 25360, 26435, 27224, 27403, 26842, 26263, 25724, 
    24925, 24283,
  25356, 25403, 26732, 26590, 26071, 25021, 23756, 23014, 22691, 22729, 
    22935, 23406, 24247, 25509, 26207, 27057, 27279, 26776, 26256, 25687, 
    24957, 24310,
  23883, 24001, 25773, 25993, 25788, 24965, 23711, 23056, 22720, 22781, 
    22993, 23473, 24267, 25703, 26195, 26187, 27060, 26784, 26221, 25756, 
    24970, 24257,
  22120, 22315, 23993, 24911, 25456, 24830, 23725, 23056, 22750, 22719, 
    22913, 23448, 24294, 25444, 26718, 24130, 25798, 26662, 26297, 25818, 
    25104, 24431,
  20668, 20908, 22617, 24227, 25167, 24732, 23677, 23012, 22770, 22788, 
    22908, 23387, 24378, 25717, 26667, 22166, 25002, 26590, 26291, 25893, 
    25193, 24471,
  20206, 20419, 22417, 24109, 25122, 24763, 23649, 23025, 22726, 22765, 
    22942, 23463, 24374, 25512, 26573, 21509, 24847, 26575, 26332, 25825, 
    25244, 24612,
  20994, 21082, 23591, 24755, 25302, 24761, 23639, 23031, 22774, 22739, 
    23008, 23446, 24293, 25536, 26689, 22650, 25090, 26597, 26346, 25893, 
    25200, 24586,
  22609, 22524, 25502, 25901, 25707, 24778, 23601, 23025, 22733, 22708, 
    22894, 23454, 24248, 25629, 26667, 25347, 26819, 26792, 26340, 25825, 
    25194, 24566,
  24203, 24013, 26740, 26467, 25851, 24820, 23594, 22963, 22751, 22803, 
    23031, 23467, 24330, 25618, 26551, 27000, 27535, 26850, 26375, 25769, 
    25258, 24613,
  25077, 24914, 26751, 26481, 25863, 24756, 23525, 22949, 22766, 22841, 
    23023, 23459, 24404, 25375, 26854, 27120, 27310, 26785, 26347, 25788, 
    25207, 24647,
  25062, 25007, 26451, 26247, 25749, 24686, 23519, 22984, 22736, 22869, 
    22997, 23510, 24510, 25541, 26418, 26876, 27235, 26676, 26251, 25795, 
    25150, 24540,
  24443, 24478, 26096, 26029, 25626, 24616, 23470, 22976, 22758, 22827, 
    23063, 23518, 24535, 25706, 26844, 26615, 27187, 26626, 26196, 25670, 
    25029, 24534,
  23610, 23680, 25774, 25907, 25563, 24526, 23432, 22949, 22752, 22816, 
    23046, 23516, 24523, 25682, 26924, 26307, 27056, 26584, 26147, 25684, 
    25030, 24494,
  22816, 22898, 25462, 25641, 25394, 24507, 23408, 22965, 22726, 22790, 
    22967, 23564, 24516, 25609, 26879, 25810, 26919, 26554, 26057, 25628, 
    24922, 24280,
  22171, 22285, 24720, 25324, 25248, 24415, 23384, 22926, 22711, 22868, 
    23055, 23493, 24543, 25756, 26837, 24692, 26490, 26534, 26057, 25616, 
    24941, 24434,
  21745, 21910, 24064, 24982, 25154, 24406, 23381, 22912, 22779, 22900, 
    23025, 23590, 24590, 25742, 27246, 23379, 25695, 26440, 26128, 25610, 
    24961, 24381,
  21584, 21775, 24175, 25028, 25132, 24342, 23350, 22939, 22756, 22843, 
    23107, 23601, 24484, 25735, 26818, 23108, 25900, 26368, 26114, 25635, 
    24961, 24495,
  21617, 21765, 24675, 25233, 25152, 24233, 23284, 22901, 22759, 22895, 
    23122, 23646, 24650, 26076, 26859, 23668, 26031, 26440, 26121, 25709, 
    25070, 24382,
  21602, 21641, 24923, 25313, 25138, 24220, 23228, 22880, 22762, 22883, 
    23102, 23646, 24662, 25889, 26882, 23787, 26062, 26498, 26107, 25784, 
    25134, 24683,
  21234, 21172, 25025, 25333, 25101, 24194, 23198, 22869, 22748, 22895, 
    23148, 23660, 24601, 25922, 26478, 23761, 26137, 26470, 26073, 25660, 
    25077, 24436,
  20432, 20335, 24893, 25308, 25061, 24161, 23177, 22834, 22751, 22921, 
    23106, 23705, 24759, 25947, 26959, 23672, 26229, 26412, 26094, 25648, 
    25032, 24423,
  19536, 19393, 24625, 25204, 24978, 24016, 23132, 22831, 22783, 22947, 
    23160, 23767, 24542, 25913, 27039, 23074, 26324, 26369, 26026, 25568, 
    25032, 24510,
  19044, 18708, 24483, 25094, 24930, 24002, 23105, 22826, 22749, 22881, 
    23095, 23729, 24658, 26079, 27247, 22379, 26193, 26326, 25978, 25450, 
    24842, 24236,
  19049, 18413, 24546, 25166, 24884, 23966, 23021, 22849, 22743, 22991, 
    23109, 23678, 24733, 26274, 27116, 22189, 26100, 26290, 25812, 25245, 
    24594, 23942,
  19145, 18356, 24739, 25204, 24827, 23837, 22987, 22761, 22755, 22879, 
    23129, 23760, 24859, 26239, 26993, 22192, 25839, 25735, 25344, 24842, 
    24130, 23608,
  28649, 28642, 27774, 27068, 25753, 24130, 22679, 22195, 22146, 22489, 
    22951, 23581, 24662, 25851, 26526, 28503, 28704, 27900, 27401, 26795, 
    25954, 25036,
  28608, 28608, 27797, 27138, 25890, 24237, 22727, 22185, 22099, 22481, 
    22818, 23581, 24607, 25522, 26570, 28503, 28729, 27893, 27353, 26775, 
    25909, 25050,
  28510, 28531, 27776, 27259, 25976, 24371, 22865, 22265, 22102, 22440, 
    22846, 23447, 24595, 25868, 26529, 28567, 28654, 27792, 27249, 26651, 
    25813, 24849,
  28403, 28452, 27824, 27191, 26104, 24457, 22938, 22300, 22110, 22486, 
    22817, 23530, 24481, 25526, 26285, 28379, 28549, 27699, 27179, 26620, 
    25762, 24989,
  28319, 28391, 27723, 27151, 26150, 24552, 22976, 22288, 22104, 22483, 
    22799, 23535, 24491, 25670, 26332, 28294, 28418, 27669, 27090, 26557, 
    25685, 24708,
  28272, 28347, 27731, 27229, 26160, 24628, 23097, 22352, 22109, 22411, 
    22728, 23412, 24621, 25651, 26610, 28232, 28400, 27698, 27104, 26532, 
    25653, 24821,
  28272, 28330, 27700, 27264, 26281, 24748, 23111, 22387, 22136, 22479, 
    22896, 23514, 24406, 25742, 26679, 28249, 28418, 27704, 27179, 26495, 
    25596, 24680,
  28319, 28359, 27865, 27379, 26347, 24810, 23211, 22460, 22135, 22384, 
    22907, 23539, 24401, 25644, 26485, 28403, 28543, 27712, 27021, 26390, 
    25366, 24567,
  28378, 28415, 27928, 27450, 26396, 24908, 23236, 22419, 22170, 22401, 
    22778, 23358, 24162, 25554, 26519, 28439, 28635, 27647, 26910, 26153, 
    25258, 24399,
  28393, 28444, 27907, 27460, 26501, 24947, 23273, 22495, 22141, 22407, 
    22713, 23487, 24243, 25579, 26431, 28442, 28579, 27568, 26814, 26072, 
    25035, 24158,
  28332, 28403, 27938, 27444, 26529, 25036, 23329, 22527, 22172, 22389, 
    22803, 23416, 24193, 25457, 26524, 28414, 28560, 27610, 26757, 26016, 
    25028, 24211,
  28221, 28308, 27862, 27468, 26575, 25027, 23363, 22568, 22181, 22454, 
    22687, 23447, 24174, 25281, 26368, 28339, 28560, 27654, 26903, 26128, 
    25041, 24325,
  28109, 28200, 27743, 27425, 26554, 25126, 23484, 22607, 22239, 22451, 
    22772, 23375, 24338, 25669, 26388, 28219, 28431, 27596, 26889, 26151, 
    25053, 24338,
  28022, 28095, 27704, 27401, 26501, 25131, 23443, 22606, 22189, 22351, 
    22794, 23443, 24340, 25569, 26184, 28129, 28331, 27568, 26793, 26015, 
    24989, 24257,
  27953, 27994, 27651, 27332, 26564, 25150, 23536, 22653, 22206, 22368, 
    22754, 23336, 24146, 25352, 26545, 28004, 28032, 27235, 26468, 25754, 
    24913, 24190,
  27900, 27917, 27565, 27293, 26547, 25147, 23546, 22682, 22262, 22413, 
    22685, 23351, 24289, 25480, 26189, 27915, 27895, 26882, 26129, 25468, 
    24702, 24156,
  27879, 27889, 27501, 27293, 26554, 25228, 23626, 22776, 22291, 22450, 
    22716, 23382, 24212, 25242, 26532, 27865, 27795, 26694, 26047, 25412, 
    24734, 24176,
  27899, 27905, 27579, 27338, 26598, 25234, 23632, 22755, 22346, 22389, 
    22745, 23272, 24256, 25140, 26445, 27915, 27739, 26571, 25922, 25312, 
    24695, 24169,
  27939, 27933, 27729, 27416, 26618, 25284, 23681, 22758, 22305, 22361, 
    22724, 23351, 24132, 25401, 26382, 28091, 27832, 26521, 25874, 25361, 
    24791, 24195,
  27963, 27943, 27778, 27429, 26698, 25317, 23719, 22749, 22319, 22404, 
    22753, 23338, 24083, 25214, 26454, 28076, 27820, 26470, 25888, 25392, 
    24746, 24142,
  27952, 27928, 27641, 27295, 26666, 25376, 23767, 22861, 22334, 22440, 
    22764, 23302, 24285, 25480, 26375, 27976, 27664, 26376, 25784, 25299, 
    24720, 24121,
  27912, 27889, 27499, 27263, 26606, 25334, 23799, 22828, 22357, 22383, 
    22664, 23299, 24203, 25300, 26026, 27771, 27228, 26354, 25832, 25373, 
    24675, 24174,
  27847, 27820, 27494, 27203, 26579, 25323, 23795, 22872, 22391, 22377, 
    22797, 23327, 24220, 25216, 26404, 27676, 27222, 26296, 25851, 25323, 
    24732, 24094,
  27737, 27694, 27539, 27287, 26560, 25410, 23798, 22880, 22406, 22414, 
    22749, 23375, 24146, 25176, 26343, 27765, 27185, 26354, 25818, 25416, 
    24744, 24120,
  27566, 27482, 27497, 27279, 26595, 25412, 23819, 22910, 22353, 22471, 
    22723, 23316, 24318, 25372, 26364, 27790, 27359, 26368, 25790, 25292, 
    24598, 24026,
  27352, 27203, 27257, 27104, 26551, 25392, 23885, 22921, 22443, 22339, 
    22808, 23369, 24207, 25241, 26667, 27659, 27291, 26318, 25741, 25161, 
    24597, 23953,
  27148, 26942, 27004, 26974, 26507, 25448, 23885, 22951, 22420, 22422, 
    22791, 23237, 24111, 25167, 26471, 27294, 26904, 26050, 25624, 25267, 
    24540, 23959,
  27005, 26796, 26837, 26879, 26497, 25392, 23905, 22977, 22408, 22441, 
    22822, 23257, 24022, 25192, 26460, 27088, 26754, 25942, 25582, 25104, 
    24508, 23952,
  26953, 26789, 26900, 26923, 26497, 25465, 23933, 23003, 22448, 22447, 
    22736, 23356, 24079, 25148, 26066, 27147, 26704, 25906, 25437, 25086, 
    24438, 23838,
  26973, 26852, 27160, 27015, 26554, 25454, 23915, 22989, 22504, 22435, 
    22699, 23391, 24113, 25245, 26309, 27306, 26554, 25876, 25409, 24998, 
    24425, 23818,
  27009, 26899, 27226, 27074, 26557, 25431, 23974, 22977, 22498, 22432, 
    22688, 23274, 24091, 25292, 26674, 27310, 26212, 25545, 25285, 24973, 
    24411, 23938,
  27001, 26880, 27185, 26976, 26537, 25451, 23964, 23050, 22495, 22507, 
    22795, 23267, 24122, 25257, 26379, 27172, 25845, 25422, 25216, 24986, 
    24418, 23844,
  26940, 26800, 26948, 26899, 26476, 25451, 23970, 23044, 22536, 22463, 
    22735, 23289, 24147, 25231, 26051, 27057, 26019, 25537, 25326, 24954, 
    24430, 23997,
  26858, 26700, 26844, 26812, 26394, 25425, 23970, 23062, 22515, 22489, 
    22741, 23332, 24105, 25177, 26119, 26999, 26119, 25674, 25436, 25091, 
    24557, 23977,
  26790, 26630, 26785, 26810, 26413, 25400, 24005, 23050, 22500, 22434, 
    22769, 23243, 24067, 25429, 26618, 26919, 26212, 25760, 25436, 25109, 
    24436, 23903,
  26746, 26604, 26726, 26737, 26359, 25364, 24005, 23088, 22547, 22443, 
    22775, 23294, 24100, 25175, 26329, 26832, 26224, 25789, 25429, 25097, 
    24487, 23950,
  26710, 26594, 26676, 26664, 26364, 25406, 24019, 23097, 22573, 22469, 
    22740, 23294, 24144, 25427, 26154, 26779, 26250, 25818, 25498, 25165, 
    24500, 23977,
  26656, 26560, 26719, 26660, 26267, 25352, 24012, 23070, 22579, 22431, 
    22821, 23263, 23912, 25413, 26489, 26744, 26349, 25912, 25594, 25190, 
    24550, 24037,
  26550, 26463, 26651, 26621, 26224, 25333, 24015, 23100, 22561, 22494, 
    22772, 23227, 24151, 25327, 26153, 26610, 26112, 25818, 25539, 25209, 
    24589, 24117,
  26368, 26282, 26623, 26553, 26232, 25366, 24046, 23120, 22593, 22517, 
    22883, 23260, 24015, 25168, 26141, 26396, 25938, 25803, 25525, 25159, 
    24537, 24144,
  26116, 26029, 26471, 26459, 26147, 25341, 24032, 23102, 22587, 22505, 
    22755, 23225, 24099, 25093, 26334, 26203, 25757, 25731, 25532, 25065, 
    24556, 24037,
  25842, 25755, 26369, 26394, 26115, 25355, 24015, 23084, 22578, 22442, 
    22777, 23280, 24104, 25287, 26213, 26237, 25907, 25810, 25525, 25202, 
    24607, 24123,
  25617, 25532, 26268, 26367, 26151, 25330, 23994, 23143, 22625, 22531, 
    22791, 23243, 24072, 25264, 26135, 26159, 26018, 25860, 25573, 25158, 
    24576, 24084,
  25505, 25414, 26174, 26346, 26113, 25301, 23990, 23149, 22602, 22459, 
    22774, 23258, 24104, 25052, 26315, 26062, 25751, 25746, 25553, 25221, 
    24588, 24144,
  25526, 25421, 26138, 26241, 26113, 25304, 23997, 23128, 22634, 22482, 
    22743, 23189, 24087, 25324, 26135, 25984, 25483, 25695, 25539, 25140, 
    24524, 24110,
  25656, 25535, 26253, 26340, 26135, 25310, 24046, 23158, 22634, 22488, 
    22791, 23334, 23968, 25399, 26697, 26048, 25907, 25695, 25525, 25158, 
    24569, 24103,
  25838, 25711, 26415, 26397, 26154, 25273, 24081, 23120, 22675, 22548, 
    22802, 23311, 24005, 25112, 26206, 26112, 25850, 25695, 25511, 25146, 
    24613, 24157,
  26019, 25896, 26359, 26462, 26184, 25341, 24029, 23149, 22666, 22548, 
    22917, 23321, 24030, 25287, 26245, 26101, 25826, 25846, 25560, 25177, 
    24652, 24130,
  26169, 26043, 26359, 26443, 26184, 25310, 24008, 23193, 22631, 22583, 
    22777, 23298, 24252, 25240, 26290, 26198, 25931, 25846, 25573, 25245, 
    24594, 24077,
  26267, 26119, 26435, 26524, 26190, 25357, 24053, 23123, 22684, 22594, 
    22717, 23324, 24119, 25361, 26504, 26293, 25900, 25731, 25497, 25208, 
    24620, 24157,
  26276, 26114, 26625, 26569, 26264, 25360, 24025, 23167, 22634, 22574, 
    22783, 23326, 24035, 25231, 26329, 26332, 25502, 25362, 25352, 25134, 
    24569, 24190,
  26166, 26026, 26499, 26534, 26226, 25293, 24039, 23137, 22651, 22560, 
    22840, 23242, 24141, 25326, 26443, 26268, 25047, 25132, 25152, 24978, 
    24512, 24144,
  25935, 25845, 26316, 26416, 26154, 25304, 24018, 23137, 22654, 22623, 
    22734, 23298, 24084, 25410, 26165, 26101, 25010, 25081, 25118, 24978, 
    24614, 24097,
  25607, 25556, 26098, 26235, 26129, 25321, 24008, 23188, 22684, 22549, 
    22797, 23296, 24166, 25231, 26334, 25892, 25054, 25103, 25069, 24978, 
    24518, 24070,
  25213, 25164, 25951, 26190, 26144, 25299, 24005, 23140, 22637, 22632, 
    22783, 23362, 24084, 25291, 26325, 25782, 25209, 25262, 25145, 24997, 
    24461, 24030,
  24806, 24731, 25851, 26092, 26069, 25271, 23987, 23140, 22655, 22580, 
    22806, 23248, 24097, 25257, 26456, 25685, 25851, 25644, 25380, 25015, 
    24607, 23996,
  24490, 24396, 25707, 25988, 26026, 25282, 23997, 23161, 22681, 22594, 
    22883, 23263, 24109, 25138, 26326, 25546, 26279, 25970, 25553, 25190, 
    24601, 24084,
  24418, 24337, 25550, 25990, 25995, 25265, 23970, 23105, 22640, 22603, 
    22758, 23327, 24126, 25434, 26554, 25354, 26529, 26244, 25747, 25171, 
    24525, 24057,
  24710, 24670, 25649, 26034, 26024, 25279, 23970, 23135, 22682, 22652, 
    22857, 23251, 24211, 25278, 26037, 25432, 26592, 26381, 25807, 25203, 
    24653, 24050,
  25359, 25357, 26139, 26332, 26160, 25277, 23984, 23147, 22705, 22672, 
    22866, 23375, 24285, 25331, 26351, 26079, 26910, 26446, 25843, 25246, 
    24634, 24057,
  26198, 26221, 26904, 26823, 26345, 25302, 23984, 23141, 22658, 22629, 
    22818, 23362, 24095, 25236, 26160, 27078, 27446, 26634, 25892, 25302, 
    24583, 24118,
  26989, 27035, 27351, 27132, 26439, 25378, 23932, 23150, 22661, 22664, 
    22775, 23309, 24137, 25373, 26201, 27651, 27576, 26713, 25982, 25377, 
    24704, 24145,
  27544, 27629, 27499, 27179, 26471, 25386, 23936, 23156, 22729, 22613, 
    22830, 23398, 24203, 25264, 26460, 27679, 27688, 26764, 26051, 25321, 
    24672, 24152,
  27811, 27945, 27453, 27154, 26432, 25330, 23911, 23144, 22717, 22679, 
    22904, 23365, 24228, 25362, 26494, 27612, 27589, 26873, 26154, 25427, 
    24736, 24306,
  27862, 28025, 27401, 27147, 26488, 25336, 23867, 23162, 22706, 22624, 
    22869, 23394, 24209, 25472, 26618, 27651, 27601, 26938, 26189, 25477, 
    24800, 24259,
  27801, 27950, 27316, 27074, 26448, 25269, 23891, 23148, 22723, 22667, 
    22929, 23381, 24177, 25236, 26441, 27620, 27732, 26923, 26210, 25514, 
    24839, 24299,
  27673, 27771, 27263, 27071, 26435, 25243, 23881, 23118, 22753, 22688, 
    22938, 23391, 24224, 25383, 26270, 27504, 27589, 26901, 26203, 25564, 
    24845, 24259,
  27444, 27484, 27220, 26974, 26359, 25238, 23839, 23054, 22715, 22671, 
    23010, 23371, 24098, 25490, 26638, 27478, 27551, 26923, 26251, 25552, 
    24794, 24280,
  27062, 27071, 27238, 26966, 26256, 25193, 23846, 23071, 22692, 22688, 
    22896, 23488, 24197, 25316, 26345, 27420, 27496, 26807, 26210, 25533, 
    24846, 24213,
  26532, 26544, 27172, 26872, 26194, 25165, 23780, 23039, 22733, 22677, 
    23036, 23420, 24155, 25386, 26460, 27381, 27490, 26829, 26169, 25559, 
    24807, 24240,
  25900, 25939, 26900, 26718, 26114, 25073, 23773, 23075, 22715, 22829, 
    22897, 23417, 24244, 25307, 26619, 27226, 27471, 26823, 26197, 25584, 
    24865, 24301,
  25158, 25246, 26513, 26481, 26010, 24989, 23756, 23046, 22745, 22720, 
    22914, 23428, 24161, 25293, 26314, 26976, 27451, 26829, 26231, 25739, 
    24948, 24267,
  24195, 24354, 26135, 26269, 25925, 24992, 23767, 23096, 22678, 22729, 
    22942, 23474, 24366, 25270, 26541, 26670, 27315, 26867, 26335, 25751, 
    25044, 24422,
  22920, 23152, 25192, 25703, 25704, 24905, 23726, 23022, 22707, 22726, 
    22928, 23451, 24287, 25430, 26525, 25513, 26867, 26729, 26342, 25790, 
    25006, 24375,
  21478, 21750, 23782, 24863, 25373, 24810, 23708, 23064, 22769, 22776, 
    22986, 23393, 24265, 25489, 26520, 23417, 25379, 26607, 26335, 25896, 
    25235, 24563,
  20335, 20583, 22870, 24346, 25172, 24754, 23684, 23038, 22734, 22796, 
    22920, 23421, 24152, 25505, 26699, 22069, 24950, 26650, 26335, 25865, 
    25236, 24509,
  20039, 20187, 22733, 24269, 25155, 24771, 23657, 22999, 22746, 22762, 
    23026, 23431, 24246, 25561, 26650, 21762, 24826, 26549, 26253, 25901, 
    25192, 24490,
  20779, 20765, 23902, 24829, 25307, 24684, 23629, 22956, 22737, 22788, 
    23026, 23455, 24406, 25607, 26375, 22973, 25418, 26615, 26295, 25828, 
    25147, 24497,
  22150, 21982, 25704, 25917, 25731, 24757, 23598, 23003, 22756, 22771, 
    23058, 23549, 24241, 25771, 26423, 25570, 27010, 26801, 26316, 25822, 
    25192, 24617,
  23392, 23165, 26632, 26447, 25820, 24797, 23529, 23018, 22720, 22800, 
    23055, 23549, 24330, 25757, 26237, 26978, 27546, 26824, 26288, 25766, 
    25045, 24624,
  23909, 23750, 26341, 26229, 25710, 24696, 23497, 22992, 22750, 22794, 
    22956, 23554, 24446, 25659, 26528, 26838, 27260, 26666, 26254, 25810, 
    25103, 24658,
  23620, 23591, 25748, 25871, 25574, 24649, 23529, 22986, 22756, 22843, 
    23053, 23534, 24506, 25718, 26746, 26151, 27035, 26594, 26178, 25704, 
    25014, 24498,
  22867, 22947, 25056, 25513, 25393, 24579, 23488, 22983, 22748, 22821, 
    23056, 23550, 24513, 25650, 26847, 25435, 26706, 26535, 26144, 25660, 
    25002, 24458,
  22067, 22206, 24580, 25279, 25337, 24492, 23418, 22960, 22792, 22827, 
    23013, 23580, 24518, 25734, 26992, 24877, 26532, 26629, 26089, 25593, 
    24932, 24358,
  21465, 21631, 24260, 25072, 25234, 24464, 23384, 22955, 22777, 22839, 
    23125, 23606, 24428, 25697, 27015, 24224, 26203, 26500, 26103, 25593, 
    24939, 24365,
  21132, 21316, 23903, 24865, 25131, 24364, 23370, 22925, 22795, 22919, 
    23037, 23594, 24514, 25881, 26569, 23367, 25829, 26515, 26062, 25631, 
    24971, 24345,
  21085, 21270, 23764, 24795, 25100, 24336, 23319, 22926, 22795, 22851, 
    23034, 23639, 24573, 25735, 26606, 22637, 25556, 26428, 26069, 25600, 
    24952, 24299,
  21311, 21462, 24231, 25035, 25114, 24319, 23367, 22894, 22787, 22888, 
    23046, 23668, 24610, 25704, 26918, 22963, 25835, 26407, 26097, 25607, 
    24870, 24372,
  21680, 21757, 24818, 25296, 25186, 24280, 23326, 22923, 22761, 22880, 
    23126, 23656, 24490, 25865, 26768, 23720, 26072, 26523, 26131, 25675, 
    25080, 24493,
  21904, 21888, 25062, 25390, 25132, 24213, 23236, 22856, 22814, 22834, 
    23137, 23587, 24473, 25870, 26899, 23949, 26160, 26435, 26090, 25650, 
    25131, 24494,
  21676, 21598, 25136, 25431, 25069, 24183, 23212, 22868, 22802, 22837, 
    23072, 23610, 24756, 25954, 26773, 24024, 26141, 26415, 26007, 25694, 
    25004, 24440,
  20933, 20846, 25088, 25380, 25049, 24124, 23195, 22859, 22785, 22938, 
    23058, 23687, 24592, 25896, 27049, 23978, 26253, 26422, 26015, 25595, 
    24954, 24380,
  20007, 19881, 24695, 25213, 24960, 24048, 23112, 22806, 22759, 22861, 
    23073, 23770, 24693, 26029, 26938, 23216, 26341, 26387, 25946, 25533, 
    24935, 24307,
  19383, 19062, 24500, 25144, 24900, 23984, 23115, 22830, 22751, 22936, 
    23102, 23768, 24782, 26159, 26609, 22276, 26129, 26285, 25891, 25403, 
    24865, 24301,
  19212, 18587, 24685, 25176, 24875, 23923, 23070, 22828, 22792, 22870, 
    23187, 23707, 24819, 25987, 27156, 22314, 26154, 26250, 25843, 25279, 
    24611, 23980,
  19224, 18445, 24941, 25251, 24801, 23800, 22981, 22769, 22772, 22893, 
    23105, 23715, 24844, 26218, 26660, 22378, 26004, 26012, 25513, 25037, 
    24288, 23573,
  28678, 28645, 27760, 27041, 25762, 24142, 22645, 22199, 22103, 22393, 
    22861, 23608, 24595, 25719, 26420, 28520, 28726, 27876, 27397, 26860, 
    25912, 24921,
  28638, 28611, 27837, 27068, 25839, 24226, 22766, 22210, 22074, 22479, 
    22860, 23562, 24644, 25604, 26335, 28498, 28769, 27920, 27363, 26625, 
    25823, 24847,
  28540, 28534, 27853, 27138, 25967, 24357, 22776, 22180, 22062, 22427, 
    22854, 23524, 24557, 25751, 26548, 28568, 28757, 27804, 27307, 26668, 
    25791, 24813,
  28429, 28461, 27728, 27197, 26060, 24438, 22883, 22242, 22067, 22473, 
    22868, 23503, 24404, 25453, 26468, 28406, 28526, 27667, 27135, 26568, 
    25726, 24826,
  28338, 28410, 27670, 27151, 26107, 24559, 22987, 22309, 22079, 22433, 
    22911, 23549, 24418, 25749, 26403, 28294, 28421, 27609, 27038, 26395, 
    25567, 24605,
  28280, 28372, 27713, 27216, 26157, 24614, 23057, 22341, 22110, 22493, 
    22760, 23483, 24546, 25667, 26823, 28174, 28359, 27674, 27093, 26394, 
    25529, 24485,
  28266, 28348, 27753, 27232, 26232, 24656, 23087, 22341, 22119, 22478, 
    22876, 23460, 24413, 25509, 26446, 28241, 28401, 27725, 27073, 26320, 
    25491, 24578,
  28298, 28353, 27812, 27320, 26344, 24768, 23157, 22406, 22098, 22446, 
    22793, 23394, 24233, 25564, 26340, 28347, 28501, 27667, 26954, 26257, 
    25280, 24410,
  28346, 28381, 27932, 27412, 26393, 24863, 23191, 22458, 22101, 22380, 
    22796, 23378, 24364, 25574, 26654, 28442, 28607, 27651, 26920, 26139, 
    25140, 24236,
  28356, 28388, 27960, 27493, 26501, 24880, 23257, 22508, 22109, 22411, 
    22812, 23507, 24550, 25625, 26529, 28487, 28670, 27645, 26893, 26070, 
    25031, 24196,
  28293, 28333, 27948, 27487, 26473, 24972, 23368, 22534, 22167, 22365, 
    22701, 23459, 24193, 25524, 26426, 28445, 28651, 27651, 26885, 26138, 
    25101, 24149,
  28179, 28230, 27847, 27450, 26544, 25022, 23389, 22561, 22179, 22425, 
    22781, 23357, 24323, 25545, 26243, 28325, 28539, 27601, 26816, 26095, 
    25063, 24135,
  28069, 28125, 27774, 27366, 26535, 25106, 23409, 22611, 22220, 22419, 
    22735, 23375, 24264, 25494, 26187, 28210, 28389, 27457, 26775, 25939, 
    24980, 24081,
  27995, 28036, 27662, 27350, 26521, 25153, 23471, 22595, 22214, 22399, 
    22786, 23435, 24281, 25442, 26732, 28079, 28234, 27284, 26504, 25815, 
    24980, 24261,
  27949, 27956, 27585, 27301, 26518, 25120, 23506, 22651, 22263, 22389, 
    22808, 23358, 24310, 25212, 26187, 27985, 27897, 26995, 26222, 25566, 
    24706, 24101,
  27915, 27892, 27563, 27266, 26515, 25136, 23551, 22662, 22301, 22406, 
    22740, 23338, 24288, 25431, 26182, 27860, 27685, 26540, 25876, 25361, 
    24705, 23993,
  27892, 27865, 27507, 27235, 26460, 25167, 23599, 22692, 22274, 22401, 
    22779, 23391, 24145, 25582, 26385, 27737, 27113, 26151, 25670, 25242, 
    24584, 24174,
  27888, 27870, 27525, 27235, 26515, 25248, 23616, 22745, 22309, 22403, 
    22756, 23345, 24216, 25344, 26226, 27659, 26939, 26078, 25656, 25192, 
    24596, 24100,
  27892, 27877, 27635, 27298, 26575, 25259, 23644, 22797, 22300, 22403, 
    22730, 23236, 24248, 25311, 26691, 27771, 26757, 26129, 25676, 25285, 
    24691, 24113,
  27882, 27863, 27540, 27368, 26606, 25293, 23706, 22812, 22344, 22411, 
    22764, 23281, 24250, 25393, 26399, 27810, 27050, 26244, 25746, 25353, 
    24729, 24079,
  27855, 27826, 27535, 27325, 26579, 25349, 23775, 22811, 22322, 22428, 
    22753, 23372, 24348, 25437, 26442, 27779, 27244, 26301, 25787, 25260, 
    24659, 24086,
  27820, 27773, 27451, 27231, 26603, 25329, 23782, 22867, 22337, 22422, 
    22701, 23316, 24237, 25311, 26485, 27659, 27362, 26279, 25710, 25204, 
    24570, 24032,
  27761, 27695, 27466, 27244, 26574, 25314, 23789, 22935, 22401, 22396, 
    22747, 23420, 24138, 25292, 26384, 27712, 27299, 26294, 25807, 25241, 
    24614, 24078,
  27645, 27569, 27471, 27293, 26576, 25390, 23803, 22875, 22348, 22399, 
    22780, 23300, 24126, 25245, 26234, 27821, 27337, 26307, 25724, 25290, 
    24639, 24011,
  27470, 27384, 27350, 27169, 26554, 25384, 23862, 22896, 22427, 22378, 
    22706, 23300, 24227, 25327, 26504, 27754, 27417, 26272, 25717, 25272, 
    24493, 24037,
  27288, 27171, 27082, 26999, 26488, 25384, 23896, 22902, 22418, 22447, 
    22740, 23320, 24096, 25141, 26335, 27515, 27293, 26250, 25703, 25228, 
    24639, 23937,
  27158, 27007, 27007, 26899, 26491, 25440, 23854, 23002, 22432, 22398, 
    22717, 23386, 24222, 25289, 26195, 27317, 27025, 25982, 25537, 25122, 
    24485, 23883,
  27100, 26955, 26996, 26894, 26528, 25389, 23875, 22984, 22441, 22515, 
    22717, 23267, 24135, 25471, 26318, 27322, 26801, 25831, 25364, 24991, 
    24460, 23876,
  27096, 27001, 27215, 27001, 26531, 25401, 23909, 22954, 22438, 22412, 
    22700, 23330, 24088, 25268, 26296, 27387, 26763, 25779, 25406, 25016, 
    24434, 23922,
  27108, 27057, 27240, 27079, 26562, 25389, 23923, 23010, 22499, 22486, 
    22771, 23261, 24152, 25364, 26473, 27389, 26639, 25694, 25357, 24978, 
    24415, 23869,
  27092, 27045, 27118, 27031, 26496, 25426, 23899, 23016, 22505, 22466, 
    22773, 23291, 24115, 25231, 26284, 27269, 26376, 25707, 25364, 24990, 
    24383, 23976,
  27015, 26945, 26971, 26845, 26428, 25426, 23972, 22998, 22502, 22462, 
    22784, 23266, 24159, 25105, 25942, 26999, 26215, 25664, 25329, 25003, 
    24408, 23935,
  26884, 26794, 26865, 26782, 26388, 25403, 23996, 23042, 22510, 22485, 
    22844, 23312, 24203, 25273, 26434, 26794, 26226, 25729, 25412, 25033, 
    24401, 23968,
  26744, 26648, 26763, 26659, 26329, 25316, 23961, 23063, 22528, 22508, 
    22696, 23281, 24129, 25210, 26519, 26682, 26172, 25779, 25467, 25083, 
    24458, 23868,
  26637, 26549, 26719, 26632, 26279, 25378, 23999, 23107, 22569, 22499, 
    22764, 23329, 24072, 25368, 26395, 26621, 25954, 25743, 25487, 25120, 
    24503, 24042,
  26577, 26500, 26743, 26621, 26218, 25302, 23999, 23074, 22586, 22545, 
    22801, 23245, 24094, 25321, 26210, 26618, 25904, 25707, 25459, 25114, 
    24541, 24015,
  26542, 26471, 26717, 26624, 26253, 25344, 23985, 23101, 22565, 22456, 
    22696, 23229, 23998, 25230, 26254, 26562, 25960, 25772, 25467, 25089, 
    24573, 24041,
  26486, 26421, 26628, 26540, 26181, 25293, 23954, 23127, 22580, 22482, 
    22781, 23280, 24082, 25272, 26157, 26498, 25941, 25735, 25418, 25039, 
    24566, 23981,
  26355, 26301, 26550, 26513, 26164, 25291, 23998, 23115, 22594, 22522, 
    22741, 23300, 24018, 25288, 26506, 26374, 25891, 25649, 25390, 25026, 
    24515, 23927,
  26122, 26078, 26412, 26467, 26118, 25318, 24026, 23091, 22553, 22533, 
    22792, 23219, 24141, 25237, 26012, 26170, 25810, 25671, 25418, 25070, 
    24483, 23954,
  25805, 25761, 26288, 26307, 26118, 25324, 23981, 23171, 22574, 22579, 
    22775, 23404, 24266, 25454, 26573, 26078, 25648, 25707, 25459, 25157, 
    24502, 24041,
  25465, 25414, 26265, 26314, 26060, 25304, 24030, 23150, 22591, 22530, 
    22800, 23280, 24131, 25342, 26187, 26028, 25779, 25772, 25494, 25157, 
    24585, 24088,
  25180, 25119, 26207, 26326, 26057, 25265, 24019, 23132, 22629, 22547, 
    22712, 23244, 24089, 25244, 26191, 25950, 25660, 25735, 25521, 25194, 
    24560, 24075,
  25022, 24939, 26194, 26270, 26032, 25276, 24016, 23177, 22588, 22562, 
    22826, 23351, 24197, 25503, 26489, 25910, 25349, 25591, 25480, 25163, 
    24521, 23980,
  25017, 24899, 26042, 26184, 26075, 25299, 24040, 23150, 22621, 22559, 
    22815, 23328, 24133, 25202, 26237, 25887, 25598, 25656, 25431, 25120, 
    24604, 23954,
  25139, 24987, 26062, 26207, 26032, 25271, 24009, 23153, 22644, 22573, 
    22780, 23303, 24232, 25132, 26357, 25864, 25579, 25497, 25335, 25026, 
    24508, 24021,
  25325, 25164, 26106, 26232, 26015, 25260, 23977, 23144, 22632, 22559, 
    22763, 23303, 24143, 25113, 26235, 25887, 25617, 25555, 25362, 25157, 
    24630, 23987,
  25522, 25376, 26116, 26306, 26089, 25318, 23974, 23153, 22620, 22539, 
    22803, 23257, 24076, 25209, 26390, 25903, 25629, 25656, 25507, 25175, 
    24649, 24081,
  25701, 25559, 26192, 26340, 26141, 25310, 24012, 23147, 22641, 22532, 
    22803, 23295, 24284, 25258, 26070, 25984, 25679, 25634, 25445, 25175, 
    24591, 24215,
  25830, 25660, 26260, 26338, 26149, 25315, 24023, 23159, 22661, 22527, 
    22806, 23292, 23982, 25144, 26247, 26056, 25760, 25642, 25493, 25244, 
    24591, 24155,
  25856, 25654, 26293, 26401, 26181, 25327, 24057, 23147, 22641, 22599, 
    22803, 23391, 23992, 25423, 26097, 26131, 25660, 25562, 25411, 25120, 
    24604, 24128,
  25735, 25536, 26248, 26365, 26141, 25315, 23984, 23171, 22720, 22527, 
    22843, 23292, 24220, 25004, 26019, 26112, 25486, 25411, 25355, 25219, 
    24610, 24094,
  25461, 25300, 26057, 26249, 26085, 25279, 23984, 23141, 22714, 22536, 
    22843, 23249, 24091, 25146, 26170, 25872, 25442, 25469, 25355, 25082, 
    24521, 24041,
  25073, 24945, 25834, 26120, 26032, 25251, 24044, 23129, 22644, 22596, 
    22794, 23287, 24091, 25398, 26584, 25585, 25610, 25497, 25293, 25088, 
    24560, 24047,
  24628, 24505, 25641, 26044, 26001, 25245, 23984, 23144, 22679, 22567, 
    22829, 23234, 24044, 25361, 26545, 25494, 25809, 25570, 25383, 25014, 
    24585, 24014,
  24191, 24055, 25595, 25960, 26001, 25254, 23978, 23112, 22697, 22556, 
    22900, 23348, 24187, 25347, 26368, 25413, 26021, 25685, 25397, 25157, 
    24636, 24054,
  23861, 23725, 25436, 25894, 25972, 25226, 23978, 23144, 22667, 22634, 
    22860, 23389, 24143, 25270, 26346, 25351, 26407, 26110, 25583, 25175, 
    24534, 24068,
  23781, 23674, 25401, 25907, 25957, 25274, 24002, 23147, 22638, 22628, 
    22880, 23359, 24188, 25246, 26274, 25290, 26613, 26270, 25722, 25232, 
    24560, 24082,
  24077, 24021, 25443, 25920, 25967, 25243, 23978, 23162, 22683, 22617, 
    22880, 23240, 24257, 25349, 26581, 25253, 26601, 26350, 25763, 25276, 
    24623, 24162,
  24767, 24752, 25771, 26066, 26035, 25274, 23981, 23115, 22653, 22694, 
    22747, 23407, 24200, 25251, 26259, 25579, 26532, 26422, 25867, 25269, 
    24675, 24055,
  25706, 25703, 26471, 26529, 26216, 25271, 23933, 23145, 22686, 22671, 
    22767, 23397, 24173, 25090, 26315, 26507, 27093, 26610, 25957, 25332, 
    24637, 24142,
  26643, 26642, 27189, 27007, 26432, 25313, 23912, 23119, 22706, 22646, 
    22844, 23336, 24233, 25279, 26376, 27401, 27579, 26740, 26032, 25407, 
    24739, 24149,
  27350, 27370, 27349, 27109, 26422, 25342, 23954, 23178, 22712, 22706, 
    22884, 23367, 24274, 25205, 26426, 27632, 27660, 26899, 26185, 25506, 
    24790, 24183,
  27722, 27788, 27420, 27112, 26451, 25280, 23892, 23101, 22751, 22612, 
    22887, 23347, 24280, 25468, 26366, 27618, 27679, 26935, 26275, 25606, 
    24815, 24330,
  27793, 27896, 27321, 27068, 26388, 25291, 23919, 23075, 22665, 22747, 
    22918, 23395, 24262, 25461, 26417, 27563, 27673, 26964, 26310, 25593, 
    24873, 24337,
  27659, 27754, 27275, 27051, 26401, 25224, 23871, 23102, 22698, 22663, 
    22941, 23360, 24162, 25466, 26528, 27582, 27585, 26921, 26241, 25587, 
    24797, 24277,
  27373, 27411, 27240, 26982, 26328, 25277, 23909, 23108, 22687, 22744, 
    22976, 23411, 24307, 25403, 26381, 27501, 27523, 26892, 26254, 25613, 
    24822, 24257,
  26911, 26881, 27238, 26918, 26285, 25219, 23875, 23093, 22693, 22721, 
    22908, 23452, 24281, 25247, 26618, 27473, 27498, 26871, 26275, 25538, 
    24823, 24344,
  26225, 26173, 27126, 26872, 26256, 25146, 23847, 23099, 22722, 22741, 
    22913, 23414, 24120, 25524, 26490, 27445, 27573, 26914, 26324, 25644, 
    24874, 24271,
  25348, 25337, 26728, 26619, 26159, 25098, 23806, 23090, 22728, 22770, 
    22885, 23394, 24197, 25420, 26565, 27260, 27542, 26856, 26296, 25713, 
    24893, 24171,
  24409, 24479, 26031, 26179, 25935, 25025, 23778, 23076, 22769, 22774, 
    22936, 23374, 24251, 25224, 26475, 26653, 27379, 26784, 26282, 25707, 
    25021, 24312,
  23525, 23677, 25252, 25725, 25735, 24947, 23750, 23064, 22737, 22751, 
    22954, 23453, 24259, 25467, 26710, 25807, 26919, 26828, 26345, 25825, 
    25072, 24339,
  22681, 22899, 24928, 25539, 25641, 24950, 23764, 23056, 22758, 22800, 
    22948, 23387, 24321, 25539, 26276, 25402, 26776, 26776, 26325, 25800, 
    25136, 24560,
  21772, 22032, 24768, 25407, 25559, 24888, 23730, 23050, 22737, 22757, 
    22912, 23458, 24351, 25513, 26918, 24891, 26651, 26776, 26387, 25931, 
    25244, 24480,
  20806, 21069, 24358, 25170, 25473, 24827, 23734, 23059, 22779, 22789, 
    22986, 23517, 24489, 25509, 26810, 23913, 25774, 26698, 26387, 25919, 
    25245, 24607,
  20049, 20256, 23967, 24931, 25373, 24785, 23678, 23024, 22753, 22806, 
    22989, 23443, 24311, 25514, 26539, 23266, 25985, 26713, 26407, 26000, 
    25168, 24655,
  19881, 19968, 23374, 24608, 25233, 24721, 23671, 23048, 22753, 22830, 
    23020, 23479, 24400, 25574, 26782, 22550, 25171, 26619, 26346, 25944, 
    25181, 24581,
  20438, 20382, 23785, 24880, 25318, 24696, 23609, 23042, 22794, 22844, 
    23038, 23436, 24398, 25521, 26551, 23204, 25588, 26656, 26332, 25863, 
    25182, 24575,
  21406, 21248, 25435, 25793, 25607, 24783, 23567, 22972, 22774, 22844, 
    23058, 23495, 24376, 25577, 26632, 25450, 26957, 26785, 26339, 25863, 
    25208, 24535,
  22191, 22029, 26034, 26103, 25707, 24766, 23568, 22995, 22833, 22825, 
    23038, 23581, 24453, 25528, 26385, 26568, 27356, 26785, 26284, 25820, 
    25106, 24555,
  22357, 22284, 25400, 25728, 25537, 24638, 23527, 23013, 22769, 22839, 
    22953, 23480, 24332, 25500, 26544, 25923, 27045, 26699, 26215, 25771, 
    25151, 24576,
  21909, 21955, 24417, 25198, 25328, 24576, 23541, 22990, 22763, 22848, 
    22925, 23485, 24372, 25606, 27171, 24727, 26310, 26562, 26168, 25671, 
    25030, 24516,
  21203, 21338, 23773, 24819, 25159, 24515, 23482, 22976, 22804, 22843, 
    23022, 23600, 24347, 25438, 26351, 23714, 25763, 26519, 26140, 25684, 
    25018, 24603,
  20626, 20802, 23472, 24695, 25125, 24459, 23444, 22985, 22752, 22897, 
    23045, 23557, 24476, 25787, 26576, 23184, 25552, 26454, 26106, 25715, 
    25043, 24443,
  20365, 20545, 23353, 24628, 25079, 24459, 23385, 22905, 22764, 22886, 
    23026, 23585, 24449, 25816, 26917, 22835, 25515, 26404, 26064, 25641, 
    24980, 24423,
  20424, 20581, 23490, 24663, 25045, 24414, 23347, 22923, 22805, 22795, 
    23054, 23565, 24550, 25895, 26806, 22603, 25484, 26368, 26113, 25635, 
    24961, 24403,
  20759, 20869, 23857, 24871, 25097, 24387, 23326, 22897, 22820, 22852, 
    23017, 23649, 24570, 25804, 27026, 22586, 25626, 26419, 26038, 25654, 
    24904, 24397,
  21312, 21360, 24428, 25073, 25148, 24351, 23313, 22941, 22805, 22924, 
    23072, 23636, 24659, 25790, 26968, 23177, 25851, 26390, 26051, 25685, 
    25006, 24544,
  21923, 21917, 24955, 25315, 25154, 24236, 23289, 22898, 22788, 22956, 
    23169, 23736, 24462, 25874, 26676, 23818, 26038, 26376, 26085, 25660, 
    24994, 24558,
  22295, 22262, 25201, 25439, 25163, 24191, 23254, 22898, 22803, 22996, 
    23078, 23660, 24712, 25795, 26975, 24032, 26088, 26398, 26072, 25748, 
    25147, 24451,
  22143, 22115, 25282, 25455, 25138, 24166, 23248, 22913, 22797, 22908, 
    23189, 23612, 24702, 25895, 26891, 24210, 26119, 26384, 26032, 25704, 
    25065, 24492,
  21435, 21429, 25166, 25466, 25109, 24133, 23213, 22866, 22845, 22922, 
    23093, 23732, 24766, 25842, 26922, 24198, 26256, 26420, 25997, 25606, 
    24855, 24432,
  20494, 20443, 24799, 25294, 24995, 24057, 23158, 22884, 22807, 22960, 
    23176, 23658, 24658, 25929, 27043, 23378, 26343, 26341, 26025, 25538, 
    24855, 24359,
  19772, 19509, 24591, 25190, 24915, 23996, 23081, 22852, 22787, 22958, 
    23179, 23826, 24991, 26238, 26835, 22465, 26095, 26312, 25846, 25383, 
    24817, 24252,
  19456, 18881, 24883, 25233, 24881, 23890, 23030, 22820, 22801, 22989, 
    23261, 23788, 24710, 26224, 27056, 22587, 26188, 26176, 25832, 25352, 
    24671, 24145,
  19396, 18666, 25075, 25332, 24821, 23826, 22975, 22793, 22799, 22964, 
    23193, 23765, 24888, 26182, 26785, 22830, 26064, 26060, 25578, 25061, 
    24347, 23758,
  28692, 28667, 27824, 27085, 25762, 24103, 22658, 22184, 22053, 22459, 
    22916, 23554, 24568, 25654, 26904, 28557, 28760, 27906, 27335, 26665, 
    25721, 24692,
  28651, 28629, 27920, 27169, 25894, 24294, 22824, 22240, 22128, 22522, 
    22859, 23585, 24630, 25897, 26899, 28539, 28824, 27798, 27267, 26576, 
    25696, 24565,
  28553, 28545, 27901, 27223, 25996, 24361, 22855, 22243, 22101, 22488, 
    22796, 23541, 24612, 25682, 26735, 28542, 28760, 27747, 27163, 26557, 
    25638, 24671,
  28443, 28473, 27862, 27234, 26039, 24464, 22900, 22287, 22115, 22450, 
    22859, 23521, 24360, 25768, 26831, 28454, 28593, 27610, 27025, 26546, 
    25663, 24638,
  28351, 28430, 27816, 27191, 26101, 24584, 22973, 22334, 22109, 22461, 
    22807, 23465, 24355, 25751, 26921, 28315, 28506, 27574, 26976, 26440, 
    25555, 24677,
  28285, 28394, 27697, 27235, 26199, 24626, 23062, 22401, 22147, 22461, 
    22909, 23462, 24554, 25860, 26515, 28206, 28394, 27551, 26970, 26334, 
    25408, 24483,
  28253, 28357, 27737, 27247, 26201, 24710, 23118, 22380, 22156, 22418, 
    22803, 23555, 24352, 25628, 26616, 28206, 28425, 27646, 26949, 26260, 
    25312, 24382,
  28259, 28333, 27791, 27341, 26316, 24791, 23197, 22448, 22135, 22437, 
    22860, 23444, 24334, 25770, 26632, 28293, 28487, 27567, 26921, 26147, 
    25070, 24194,
  28284, 28331, 27957, 27454, 26396, 24864, 23242, 22465, 22144, 22483, 
    22829, 23522, 24329, 25584, 26279, 28393, 28606, 27631, 26859, 26048, 
    25051, 24154,
  28284, 28319, 27982, 27489, 26482, 24922, 23363, 22542, 22161, 22494, 
    22820, 23359, 24374, 25462, 26760, 28469, 28674, 27624, 26804, 26016, 
    24942, 24147,
  28226, 28261, 27973, 27500, 26484, 25034, 23349, 22556, 22184, 22453, 
    22757, 23392, 24304, 25462, 26509, 28416, 28606, 27581, 26776, 26054, 
    24923, 24046,
  28125, 28160, 27915, 27454, 26542, 25045, 23398, 22594, 22207, 22413, 
    22820, 23361, 24376, 25304, 26907, 28301, 28493, 27529, 26748, 25929, 
    24955, 24166,
  28028, 28054, 27813, 27403, 26604, 25073, 23470, 22650, 22242, 22381, 
    22785, 23379, 24333, 25546, 26382, 28126, 28344, 27292, 26589, 25779, 
    24942, 24112,
  27968, 27969, 27696, 27326, 26481, 25129, 23547, 22694, 22277, 22470, 
    22736, 23338, 24264, 25555, 26850, 28067, 28126, 27053, 26389, 25667, 
    24719, 24132,
  27937, 27906, 27618, 27295, 26524, 25132, 23504, 22693, 22247, 22381, 
    22756, 23371, 24380, 25508, 26499, 27956, 27857, 26685, 25989, 25369, 
    24648, 24012,
  27910, 27862, 27534, 27195, 26460, 25103, 23577, 22646, 22276, 22452, 
    22792, 23282, 24328, 25455, 26173, 27794, 27391, 26281, 25732, 25201, 
    24629, 24005,
  27879, 27838, 27420, 27163, 26410, 25168, 23598, 22775, 22302, 22429, 
    22781, 23350, 24219, 25438, 26281, 27467, 26768, 26007, 25601, 25139, 
    24520, 24011,
  27847, 27826, 27387, 27125, 26432, 25184, 23625, 22742, 22307, 22466, 
    22786, 23352, 24253, 25284, 26560, 27253, 25872, 25682, 25519, 25169, 
    24635, 24145,
  27813, 27807, 27460, 27168, 26524, 25218, 23684, 22804, 22310, 22425, 
    22780, 23433, 24221, 25524, 26476, 27390, 26195, 25841, 25650, 25237, 
    24602, 24178,
  27772, 27773, 27499, 27232, 26581, 25296, 23688, 22831, 22328, 22356, 
    22820, 23266, 24248, 25536, 26697, 27593, 26768, 26093, 25704, 25243, 
    24653, 24277,
  27737, 27731, 27485, 27307, 26604, 25330, 23767, 22816, 22368, 22528, 
    22728, 23341, 24169, 25268, 26225, 27632, 27310, 26279, 25760, 25237, 
    24704, 24170,
  27715, 27682, 27454, 27313, 26590, 25349, 23799, 22865, 22432, 22453, 
    22731, 23377, 24169, 25540, 26354, 27660, 27409, 26345, 25779, 25249, 
    24684, 24190,
  27673, 27612, 27503, 27300, 26554, 25358, 23809, 22874, 22423, 22450, 
    22856, 23280, 24329, 25542, 26631, 27750, 27278, 26351, 25759, 25292, 
    24633, 24002,
  27566, 27496, 27442, 27204, 26566, 25360, 23784, 22897, 22400, 22447, 
    22839, 23300, 24299, 25556, 26432, 27775, 27278, 26331, 25662, 25155, 
    24639, 24049,
  27404, 27340, 27237, 27098, 26524, 25338, 23815, 22927, 22408, 22507, 
    22759, 23320, 24326, 25197, 26348, 27575, 27216, 26207, 25635, 25056, 
    24499, 24009,
  27266, 27192, 26932, 26934, 26417, 25338, 23853, 22941, 22443, 22449, 
    22790, 23343, 24227, 25484, 26551, 27363, 26942, 25976, 25559, 25124, 
    24485, 23921,
  27209, 27119, 27031, 27017, 26476, 25371, 23895, 22968, 22440, 22489, 
    22776, 23289, 24318, 25134, 26389, 27321, 26892, 25954, 25517, 25018, 
    24447, 23927,
  27222, 27146, 27237, 27090, 26510, 25371, 23864, 22952, 22463, 22526, 
    22866, 23327, 24259, 25206, 26619, 27494, 26810, 25932, 25413, 25012, 
    24364, 23887,
  27254, 27227, 27279, 27129, 26506, 25424, 23929, 22964, 22501, 22509, 
    22792, 23314, 24027, 25414, 26429, 27535, 26767, 25846, 25399, 24980, 
    24396, 23833,
  27256, 27267, 27300, 27079, 26474, 25413, 23922, 22999, 22501, 22457, 
    22841, 23347, 24217, 25229, 26689, 27516, 26767, 25832, 25392, 25036, 
    24364, 23813,
  27200, 27200, 27173, 27022, 26449, 25379, 23950, 23038, 22509, 22437, 
    22832, 23301, 24174, 25297, 26476, 27249, 26587, 25831, 25482, 24980, 
    24459, 23880,
  27069, 27038, 26950, 26832, 26345, 25418, 23984, 23013, 22524, 22520, 
    22843, 23314, 24095, 25271, 26546, 26859, 26175, 25694, 25433, 24992, 
    24446, 24007,
  26880, 26835, 26810, 26747, 26334, 25387, 23957, 23055, 22541, 22511, 
    22868, 23326, 24196, 25371, 26185, 26585, 25690, 25528, 25371, 25048, 
    24477, 24047,
  26683, 26649, 26726, 26642, 26271, 25373, 23998, 23058, 22570, 22551, 
    22757, 23324, 24174, 25259, 26454, 26429, 25397, 25412, 25281, 25104, 
    24535, 23933,
  26530, 26513, 26751, 26564, 26257, 25322, 23967, 23122, 22541, 22525, 
    22808, 23270, 24258, 25233, 26404, 26346, 25328, 25441, 25343, 24992, 
    24426, 23973,
  26447, 26429, 26682, 26574, 26188, 25278, 23984, 23105, 22529, 22508, 
    22802, 23338, 24275, 25464, 26270, 26335, 25434, 25412, 25239, 24911, 
    24477, 23959,
  26413, 26378, 26709, 26596, 26210, 25362, 24015, 23110, 22573, 22522, 
    22817, 23316, 24124, 25084, 26444, 26313, 25639, 25571, 25350, 25010, 
    24547, 24006,
  26368, 26322, 26650, 26550, 26162, 25325, 24012, 23119, 22573, 22530, 
    22856, 23290, 24208, 25322, 26487, 26226, 25757, 25621, 25446, 25041, 
    24540, 24086,
  26241, 26207, 26524, 26509, 26147, 25314, 24005, 23125, 22623, 22487, 
    22760, 23341, 24163, 25161, 26360, 26090, 25496, 25549, 25426, 25109, 
    24598, 24066,
  25995, 25979, 26439, 26415, 26162, 25297, 23983, 23077, 22590, 22596, 
    22805, 23318, 24102, 25298, 26328, 26035, 25409, 25527, 25446, 25060, 
    24579, 24046,
  25646, 25637, 26224, 26329, 26159, 25339, 24049, 23157, 22640, 22513, 
    22785, 23338, 24252, 25240, 26560, 26007, 25770, 25671, 25467, 25072, 
    24560, 24032,
  25256, 25241, 26173, 26224, 26053, 25246, 24036, 23107, 22593, 22536, 
    22745, 23272, 24131, 25291, 26291, 25882, 25664, 25700, 25487, 25090, 
    24527, 24065,
  24906, 24881, 26082, 26194, 26064, 25291, 24015, 23172, 22616, 22550, 
    22802, 23315, 24195, 25280, 26185, 25804, 25284, 25584, 25405, 25059, 
    24496, 24045,
  24681, 24633, 25979, 26140, 26035, 25302, 24011, 23130, 22625, 22642, 
    22776, 23251, 24287, 25333, 26487, 25765, 25576, 25628, 25481, 25134, 
    24597, 23991,
  24627, 24534, 25912, 26135, 26076, 25311, 23997, 23145, 22660, 22567, 
    22804, 23315, 24202, 25261, 26003, 25723, 25614, 25570, 25383, 25134, 
    24502, 24012,
  24724, 24582, 25975, 26124, 26041, 25291, 24091, 23169, 22657, 22581, 
    22839, 23327, 24027, 25478, 26613, 25687, 25321, 25418, 25335, 25065, 
    24610, 24065,
  24905, 24740, 25957, 26143, 26053, 25291, 24029, 23166, 22710, 22598, 
    22816, 23315, 24153, 25303, 26419, 25709, 25290, 25440, 25301, 25134, 
    24648, 24139,
  25110, 24956, 26110, 26224, 26110, 25269, 24004, 23169, 22651, 22541, 
    22842, 23203, 24017, 25401, 26197, 25782, 25134, 25281, 25204, 25040, 
    24489, 24099,
  25303, 25160, 26247, 26310, 26110, 25322, 24070, 23186, 22684, 22584, 
    22830, 23343, 24116, 25158, 26323, 25943, 25396, 25368, 25287, 25028, 
    24591, 24092,
  25448, 25282, 26242, 26388, 26153, 25328, 24022, 23160, 22713, 22559, 
    22790, 23206, 24116, 25261, 26435, 26026, 25545, 25483, 25383, 25078, 
    24470, 24092,
  25486, 25278, 26191, 26321, 26104, 25347, 24018, 23145, 22684, 22544, 
    22825, 23299, 24072, 25254, 26410, 25904, 25358, 25361, 25314, 25096, 
    24546, 24052,
  25359, 25133, 26117, 26262, 26160, 25291, 24015, 23175, 22689, 22587, 
    22754, 23373, 24185, 25203, 26381, 25868, 25496, 25491, 25398, 25072, 
    24540, 24052,
  25047, 24837, 25912, 26221, 26084, 25322, 24029, 23204, 22692, 22619, 
    22862, 23333, 24163, 25196, 26510, 25760, 25913, 25714, 25494, 25140, 
    24610, 24119,
  24590, 24402, 25772, 26046, 26067, 25305, 24053, 23181, 22701, 22653, 
    22856, 23376, 24166, 25201, 26465, 25554, 26112, 25787, 25459, 25153, 
    24630, 24039,
  24065, 23888, 25613, 25971, 26018, 25249, 24067, 23175, 22681, 22565, 
    22865, 23376, 24059, 25247, 26173, 25411, 26119, 25888, 25543, 25066, 
    24508, 24153,
  23566, 23400, 25468, 25887, 25947, 25252, 24012, 23166, 22727, 22673, 
    22899, 23269, 24154, 25245, 26241, 25303, 26379, 26082, 25626, 25177, 
    24649, 24139,
  23205, 23061, 25070, 25669, 25896, 25246, 24025, 23187, 22733, 22645, 
    22788, 23356, 24205, 25424, 26403, 24988, 26435, 26199, 25709, 25215, 
    24604, 24206,
  23109, 23002, 24994, 25650, 25850, 25238, 24032, 23175, 22702, 22656, 
    22902, 23374, 24042, 25275, 26567, 24796, 26331, 26249, 25709, 25109, 
    24547, 24066,
  23390, 23325, 25156, 25720, 25881, 25264, 23953, 23134, 22678, 22657, 
    22837, 23379, 24124, 25341, 26574, 24960, 26510, 26357, 25860, 25197, 
    24585, 24093,
  24073, 24029, 25428, 25917, 25984, 25264, 23987, 23190, 22755, 22740, 
    22862, 23328, 24270, 25289, 26112, 25168, 26573, 26509, 25929, 25328, 
    24623, 24126,
  25035, 24980, 26107, 26329, 26176, 25267, 23980, 23143, 22711, 22674, 
    22919, 23369, 24085, 25483, 26270, 25971, 26798, 26726, 26082, 25452, 
    24732, 24214,
  26033, 25958, 26985, 26895, 26362, 25320, 23963, 23131, 22711, 22720, 
    22922, 23300, 24179, 25247, 26201, 27107, 27582, 26754, 26117, 25508, 
    24726, 24187,
  26816, 26751, 27404, 27067, 26449, 25292, 23936, 23111, 22731, 22680, 
    22877, 23356, 24196, 25346, 26471, 27564, 27739, 26892, 26151, 25502, 
    24777, 24234,
  27237, 27218, 27359, 27095, 26428, 25300, 23915, 23182, 22717, 22686, 
    23034, 23354, 24078, 25264, 26321, 27578, 27632, 26885, 26144, 25446, 
    24777, 24274,
  27287, 27322, 27323, 27062, 26382, 25255, 23953, 23123, 22720, 22718, 
    22969, 23346, 24155, 25374, 26047, 27504, 27582, 26864, 26235, 25583, 
    24841, 24322,
  27042, 27098, 27300, 27025, 26345, 25253, 23884, 23149, 22737, 22755, 
    22866, 23377, 24145, 25215, 26214, 27469, 27515, 26900, 26269, 25615, 
    24892, 24302,
  26570, 26598, 27212, 26981, 26310, 25222, 23915, 23123, 22776, 22753, 
    22917, 23364, 24318, 25315, 26696, 27466, 27626, 26914, 26310, 25696, 
    24969, 24315,
  25869, 25854, 26894, 26720, 26176, 25082, 23867, 23109, 22703, 22735, 
    22961, 23444, 24251, 25348, 26592, 27360, 27626, 26944, 26407, 25907, 
    25014, 24476,
  24914, 24897, 26385, 26426, 26071, 25141, 23846, 23132, 22723, 22699, 
    23003, 23474, 24276, 25250, 26570, 27045, 27646, 26915, 26366, 25839, 
    25014, 24457,
  23766, 23807, 25662, 25947, 25810, 25012, 23812, 23062, 22727, 22802, 
    22972, 23472, 24284, 25414, 26493, 26284, 27378, 26915, 26414, 25771, 
    25084, 24457,
  22615, 22740, 24445, 25250, 25524, 24939, 23798, 23091, 22751, 22782, 
    22958, 23350, 24242, 25509, 26813, 24980, 26506, 26778, 26346, 25901, 
    25104, 24578,
  21672, 21857, 23456, 24652, 25342, 24844, 23770, 23068, 22774, 22757, 
    22947, 23389, 24291, 25526, 26544, 23751, 25460, 26612, 26401, 25889, 
    25180, 24585,
  20996, 21206, 23357, 24631, 25318, 24867, 23767, 23098, 22751, 22800, 
    22973, 23374, 24447, 25533, 26676, 23528, 25411, 26648, 26374, 26001, 
    25276, 24692,
  20469, 20688, 24004, 25016, 25425, 24836, 23691, 23077, 22757, 22777, 
    22933, 23483, 24412, 25428, 26747, 24029, 25982, 26684, 26388, 25970, 
    25174, 24551,
  19970, 20186, 24841, 25420, 25579, 24932, 23764, 23104, 22775, 22855, 
    22922, 23559, 24282, 25503, 26585, 24669, 26401, 26764, 26367, 25939, 
    25238, 24672,
  19564, 19739, 24704, 25369, 25531, 24836, 23677, 23060, 22813, 22783, 
    22982, 23374, 24388, 25682, 26578, 24619, 26929, 26793, 26374, 25846, 
    25251, 24552,
  19464, 19548, 23566, 24755, 25273, 24761, 23622, 22993, 22798, 22847, 
    23013, 23456, 24293, 25591, 26576, 23192, 25754, 26569, 26291, 25859, 
    25207, 24512,
  19776, 19759, 23300, 24656, 25236, 24708, 23611, 23049, 22799, 22830, 
    22900, 23527, 24384, 25601, 26842, 22876, 25131, 26504, 26257, 25785, 
    25226, 24747,
  20307, 20240, 24423, 25224, 25411, 24714, 23632, 23022, 22764, 22888, 
    23005, 23578, 24374, 25466, 26704, 24612, 26575, 26721, 26285, 25791, 
    25227, 24633,
  20672, 20635, 24753, 25383, 25474, 24711, 23553, 23085, 22790, 22816, 
    23014, 23436, 24397, 25746, 26535, 25334, 27048, 26700, 26257, 25779, 
    25246, 24741,
  20606, 20654, 24000, 25006, 25297, 24650, 23567, 23008, 22744, 22836, 
    23020, 23464, 24333, 25592, 26765, 24321, 26140, 26554, 26189, 25742, 
    25126, 24734,
  20181, 20314, 23314, 24535, 25114, 24535, 23536, 22991, 22773, 22882, 
    23024, 23526, 24538, 25625, 26596, 23153, 25418, 26469, 26140, 25699, 
    25094, 24594,
  19724, 19901, 22883, 24377, 25063, 24513, 23491, 22962, 22827, 22857, 
    23101, 23498, 24414, 25720, 26669, 22447, 25393, 26484, 26147, 25667, 
    25075, 24541,
  19534, 19708, 22944, 24366, 25049, 24448, 23464, 23009, 22830, 22854, 
    23041, 23510, 24388, 25690, 26760, 22243, 25437, 26448, 26079, 25631, 
    25082, 24561,
  19702, 19833, 23256, 24549, 25043, 24457, 23439, 22977, 22809, 22961, 
    23107, 23483, 24499, 25639, 26884, 22279, 25550, 26426, 26093, 25704, 
    25088, 24495,
  20151, 20212, 23745, 24768, 25100, 24438, 23395, 22933, 22801, 22824, 
    23133, 23590, 24519, 25710, 26719, 22635, 25643, 26441, 25982, 25619, 
    24942, 24488,
  20790, 20773, 24303, 25021, 25140, 24368, 23370, 22936, 22739, 22941, 
    23144, 23570, 24645, 25891, 26698, 23070, 25904, 26404, 26066, 25638, 
    24949, 24509,
  21548, 21476, 24704, 25207, 25143, 24303, 23336, 22934, 22810, 22956, 
    23111, 23491, 24497, 25928, 26779, 23532, 25929, 26391, 26059, 25594, 
    25019, 24422,
  22277, 22205, 25071, 25347, 25163, 24259, 23291, 22928, 22807, 22841, 
    23057, 23669, 24546, 25728, 26717, 23861, 25973, 26434, 26128, 25650, 
    25083, 24542,
  22705, 22685, 25248, 25422, 25149, 24220, 23253, 22890, 22825, 22908, 
    23151, 23687, 24470, 25994, 27189, 24036, 25967, 26391, 26079, 25638, 
    25115, 24603,
  22581, 22633, 25289, 25482, 25084, 24175, 23267, 22896, 22773, 23005, 
    23131, 23622, 24687, 25800, 26879, 24320, 26129, 26442, 26018, 25682, 
    25020, 24630,
  21899, 21998, 25320, 25457, 25112, 24139, 23181, 22911, 22785, 22931, 
    23100, 23668, 24592, 25966, 26679, 24414, 26254, 26385, 25942, 25508, 
    24925, 24463,
  20962, 21007, 24955, 25312, 25015, 24047, 23174, 22894, 22788, 22969, 
    23237, 23784, 24762, 26003, 26684, 23552, 26266, 26392, 26053, 25607, 
    24944, 24396,
  20174, 19996, 24674, 25216, 24921, 23977, 23153, 22879, 22850, 22934, 
    23146, 23810, 24632, 26048, 26740, 22664, 26142, 26276, 25922, 25459, 
    24868, 24323,
  19743, 19257, 24975, 25318, 24887, 23904, 23112, 22862, 22818, 22969, 
    23189, 23747, 24745, 26181, 27259, 22945, 26142, 26254, 25804, 25385, 
    24760, 24196,
  19622, 18987, 25183, 25342, 24842, 23840, 23036, 22803, 22803, 22932, 
    23238, 23800, 24859, 26404, 27214, 23174, 26167, 26104, 25682, 25180, 
    24576, 23943,
  28696, 28681, 27854, 27100, 25747, 24096, 22699, 22205, 22066, 22490, 
    22757, 23521, 24667, 25771, 26722, 28624, 28782, 27884, 27318, 26638, 
    25640, 24577,
  28655, 28641, 27849, 27197, 25890, 24275, 22772, 22257, 22095, 22538, 
    22973, 23554, 24627, 25917, 26767, 28616, 28845, 27884, 27262, 26526, 
    25632, 24616,
  28559, 28556, 27918, 27282, 25967, 24379, 22868, 22245, 22127, 22515, 
    22918, 23663, 24642, 25714, 26673, 28557, 28764, 27776, 27166, 26476, 
    25557, 24529,
  28456, 28488, 27851, 27310, 26098, 24474, 22924, 22277, 22091, 22526, 
    22887, 23629, 24521, 25714, 26423, 28529, 28559, 27668, 27054, 26451, 
    25537, 24629,
  28372, 28450, 27763, 27224, 26143, 24566, 23038, 22345, 22103, 22520, 
    22935, 23629, 24404, 25672, 26765, 28385, 28422, 27567, 27054, 26438, 
    25505, 24562,
  28303, 28414, 27776, 27242, 26178, 24572, 23055, 22368, 22138, 22468, 
    22803, 23507, 24441, 25481, 26668, 28307, 28478, 27574, 26965, 26295, 
    25384, 24521,
  28250, 28362, 27750, 27257, 26232, 24745, 23104, 22409, 22146, 22468, 
    22818, 23456, 24470, 25765, 26510, 28269, 28384, 27639, 26931, 26157, 
    25155, 24320,
  28222, 28312, 27765, 27301, 26304, 24784, 23159, 22397, 22137, 22479, 
    22860, 23456, 24438, 25616, 26504, 28272, 28459, 27595, 26876, 26084, 
    25072, 24246,
  28213, 28281, 27884, 27369, 26378, 24865, 23273, 22476, 22163, 22556, 
    22814, 23491, 24364, 25450, 26474, 28473, 28571, 27674, 26985, 26090, 
    25059, 24199,
  28194, 28257, 27876, 27409, 26406, 24938, 23290, 22446, 22192, 22418, 
    22802, 23539, 24371, 25714, 26682, 28456, 28557, 27523, 26826, 25940, 
    24969, 24119,
  28138, 28200, 27879, 27393, 26482, 25016, 23352, 22555, 22224, 22449, 
    22777, 23445, 24216, 25700, 26597, 28392, 28490, 27357, 26613, 25866, 
    24912, 23991,
  28050, 28099, 27782, 27401, 26512, 25080, 23384, 22581, 22179, 22475, 
    22754, 23445, 24309, 25352, 26512, 28275, 28290, 27350, 26544, 25853, 
    24918, 24078,
  27963, 27986, 27712, 27344, 26515, 25088, 23443, 22598, 22226, 22394, 
    22742, 23432, 24319, 25536, 26481, 28160, 28166, 27104, 26412, 25598, 
    24656, 24131,
  27908, 27902, 27607, 27301, 26476, 25094, 23484, 22654, 22220, 22494, 
    22855, 23355, 24351, 25359, 26672, 27996, 27929, 26685, 25978, 25299, 
    24605, 23977,
  27881, 27854, 27613, 27250, 26454, 25147, 23515, 22610, 22252, 22442, 
    22735, 23360, 24306, 25499, 26599, 27890, 27624, 26410, 25798, 25206, 
    24567, 24063,
  27857, 27827, 27524, 27188, 26417, 25102, 23584, 22704, 22307, 22445, 
    22832, 23428, 24210, 25538, 26819, 27656, 27431, 26259, 25653, 25094, 
    24547, 24030,
  27818, 27798, 27389, 27085, 26365, 25149, 23591, 22727, 22260, 22447, 
    22832, 23340, 24323, 25359, 26739, 27382, 26807, 26021, 25570, 25125, 
    24464, 23989,
  27765, 27755, 27285, 27088, 26403, 25127, 23622, 22762, 22301, 22427, 
    22792, 23344, 24222, 25340, 26592, 27120, 25948, 25768, 25507, 25125, 
    24585, 24076,
  27702, 27699, 27429, 27153, 26501, 25219, 23694, 22777, 22327, 22479, 
    22868, 23410, 24206, 25563, 26532, 27301, 26428, 25912, 25535, 25093, 
    24552, 23988,
  27641, 27643, 27448, 27225, 26534, 25281, 23740, 22836, 22350, 22504, 
    22831, 23334, 24270, 25309, 26360, 27585, 27020, 25999, 25527, 25149, 
    24546, 24068,
  27606, 27603, 27435, 27217, 26588, 25348, 23746, 22853, 22356, 22478, 
    22820, 23356, 24159, 25437, 26591, 27631, 27219, 26135, 25685, 25173, 
    24635, 24156,
  27600, 27576, 27519, 27265, 26637, 25367, 23781, 22829, 22379, 22429, 
    22793, 23303, 24203, 25509, 26431, 27707, 27399, 26265, 25754, 25260, 
    24628, 24188,
  27576, 27531, 27597, 27290, 26594, 25373, 23836, 22885, 22387, 22517, 
    22773, 23353, 24191, 25563, 25879, 27838, 27518, 26359, 25796, 25223, 
    24602, 24128,
  27489, 27442, 27429, 27195, 26562, 25373, 23874, 22956, 22411, 22540, 
    22759, 23416, 24173, 25432, 26472, 27748, 27374, 26279, 25699, 25216, 
    24596, 24195,
  27361, 27328, 27181, 27015, 26442, 25370, 23878, 22949, 22478, 22563, 
    22722, 23378, 24311, 25299, 26566, 27470, 27137, 26142, 25541, 25067, 
    24449, 23859,
  27277, 27246, 27097, 26950, 26404, 25297, 23836, 22970, 22433, 22462, 
    22858, 23279, 24244, 25376, 26054, 27329, 26876, 25918, 25485, 25041, 
    24410, 23940,
  27284, 27247, 27237, 27054, 26490, 25358, 23863, 22975, 22500, 22531, 
    22821, 23312, 24326, 25373, 26832, 27448, 26857, 25954, 25601, 25035, 
    24448, 23765,
  27346, 27326, 27332, 27141, 26507, 25383, 23912, 22972, 22500, 22502, 
    22786, 23385, 24232, 25483, 26678, 27590, 26994, 26048, 25601, 25141, 
    24467, 23966,
  27393, 27416, 27429, 27106, 26493, 25386, 23911, 23022, 22477, 22548, 
    22855, 23359, 24089, 25373, 26397, 27621, 27081, 26106, 25629, 25134, 
    24480, 23932,
  27382, 27426, 27338, 27039, 26462, 25352, 23922, 23046, 22491, 22456, 
    22809, 23296, 24115, 25264, 26437, 27478, 26956, 26069, 25588, 25115, 
    24499, 23925,
  27297, 27315, 27166, 26904, 26407, 25372, 23960, 23016, 22514, 22533, 
    22860, 23278, 24137, 25431, 26619, 27231, 26501, 25838, 25491, 25103, 
    24524, 24012,
  27127, 27105, 26993, 26794, 26350, 25358, 23974, 23099, 22529, 22470, 
    22837, 23329, 24021, 25322, 26290, 26918, 25785, 25506, 25304, 25028, 
    24485, 24059,
  26885, 26854, 26856, 26704, 26304, 25341, 23967, 23077, 22514, 22507, 
    22780, 23359, 24145, 25375, 26159, 26651, 25230, 25087, 25145, 24891, 
    24422, 23991,
  26620, 26611, 26734, 26659, 26301, 25360, 24057, 23065, 22543, 22553, 
    22720, 23361, 24203, 25343, 26621, 26437, 25131, 25058, 25104, 24928, 
    24441, 23931,
  26400, 26409, 26635, 26582, 26212, 25299, 24012, 23080, 22549, 22607, 
    22817, 23270, 24241, 25296, 26485, 26326, 25180, 25137, 25097, 24859, 
    24389, 23998,
  26271, 26266, 26600, 26582, 26223, 25312, 24022, 23107, 22592, 22567, 
    22856, 23297, 24137, 25212, 26539, 26273, 25349, 25267, 25152, 24890, 
    24440, 23924,
  26228, 26188, 26551, 26529, 26189, 25338, 23994, 23101, 22586, 22575, 
    22796, 23226, 24198, 25247, 26493, 26203, 25330, 25310, 25193, 24921, 
    24459, 23964,
  26208, 26146, 26660, 26543, 26185, 25296, 24008, 23104, 22557, 22523, 
    22919, 23282, 23971, 25370, 26447, 26139, 25336, 25332, 25290, 24990, 
    24580, 23957,
  26126, 26072, 26645, 26462, 26192, 25332, 24018, 23162, 22604, 22517, 
    22813, 23396, 24112, 25555, 26601, 26178, 25479, 25432, 25303, 25033, 
    24542, 23977,
  25920, 25887, 26457, 26432, 26181, 25343, 24060, 23141, 22604, 22534, 
    22782, 23358, 24225, 25393, 26374, 26167, 25871, 25626, 25421, 25033, 
    24529, 24057,
  25587, 25567, 26318, 26437, 26132, 25298, 24053, 23153, 22668, 22538, 
    22896, 23401, 24161, 25253, 26029, 26067, 25846, 25728, 25434, 25064, 
    24529, 24017,
  25175, 25159, 26237, 26343, 26140, 25312, 24046, 23180, 22647, 22589, 
    22836, 23315, 24166, 25403, 25822, 25932, 25535, 25613, 25414, 25076, 
    24484, 24145,
  24773, 24753, 26104, 26204, 26103, 25298, 24035, 23165, 22656, 22560, 
    22913, 23241, 24087, 25331, 26585, 25753, 25236, 25468, 25414, 25039, 
    24491, 24057,
  24483, 24444, 25816, 26039, 25997, 25326, 24042, 23168, 22671, 22569, 
    22782, 23251, 24205, 25218, 26415, 25632, 25092, 25309, 25241, 25014, 
    24580, 24044,
  24372, 24289, 25729, 26073, 26046, 25318, 24056, 23180, 22641, 22632, 
    22952, 23413, 24195, 25284, 26404, 25577, 25036, 25338, 25324, 25101, 
    24561, 24184,
  24431, 24295, 25816, 26089, 26054, 25332, 24056, 23194, 22688, 22597, 
    22924, 23322, 24232, 25386, 26466, 25574, 25254, 25338, 25303, 25008, 
    24528, 24117,
  24596, 24428, 25831, 26073, 26063, 25320, 24035, 23209, 22720, 22574, 
    22875, 23264, 24257, 25167, 26541, 25510, 25099, 25259, 25296, 25101, 
    24624, 24198,
  24798, 24635, 25831, 26089, 26074, 25329, 24056, 23188, 22694, 22612, 
    22935, 23266, 24198, 25451, 26495, 25491, 24881, 25194, 25269, 25120, 
    24573, 24111,
  24994, 24846, 25957, 26173, 26098, 25329, 24070, 23206, 22700, 22597, 
    22901, 23357, 24141, 25191, 26497, 25716, 25329, 25446, 25358, 25039, 
    24561, 24117,
  25143, 24983, 26145, 26284, 26149, 25349, 24028, 23200, 22683, 22635, 
    22878, 23360, 24215, 25216, 26522, 25917, 25672, 25598, 25483, 25126, 
    24656, 24191,
  25187, 24990, 26128, 26319, 26146, 25326, 24098, 23224, 22683, 22637, 
    23035, 23350, 24151, 25281, 26750, 25875, 25485, 25439, 25351, 25032, 
    24554, 24164,
  25058, 24836, 26018, 26213, 26089, 25312, 24035, 23194, 22694, 22632, 
    22932, 23396, 24138, 25342, 26684, 25747, 25697, 25541, 25358, 25151, 
    24573, 24037,
  24721, 24503, 25859, 26165, 26089, 25357, 24053, 23194, 22700, 22629, 
    22910, 23345, 24262, 25325, 26541, 25638, 25853, 25591, 25310, 25120, 
    24650, 24064,
  24203, 24007, 25632, 26022, 26029, 25315, 24042, 23197, 22689, 22632, 
    22827, 23421, 24161, 25268, 26389, 25460, 26026, 25772, 25455, 25095, 
    24637, 24050,
  23596, 23427, 25418, 25904, 25931, 25295, 24053, 23192, 22724, 22663, 
    22844, 23289, 24235, 25377, 26329, 25315, 26382, 26054, 25600, 25107, 
    24567, 24191,
  23028, 22888, 24956, 25634, 25851, 25270, 24042, 23195, 22762, 22666, 
    22870, 23396, 24264, 25216, 26713, 24889, 26532, 26204, 25669, 25213, 
    24593, 24098,
  22622, 22514, 24545, 25378, 25794, 25236, 24011, 23233, 22706, 22690, 
    22887, 23381, 24225, 25519, 26376, 24271, 26151, 26364, 25787, 25170, 
    24612, 24131,
  22481, 22400, 24568, 25362, 25765, 25250, 24018, 23218, 22709, 22612, 
    22816, 23274, 24230, 25272, 26139, 24171, 26001, 26357, 25842, 25176, 
    24561, 24105,
  22680, 22609, 24845, 25532, 25837, 25234, 24005, 23177, 22706, 22652, 
    22891, 23368, 24413, 25312, 26454, 24510, 26401, 26459, 25932, 25319, 
    24657, 24105,
  23233, 23148, 25071, 25635, 25863, 25234, 23959, 23174, 22698, 22718, 
    22993, 23384, 24245, 25543, 26347, 24833, 26457, 26632, 25988, 25363, 
    24695, 24152,
  24049, 23931, 25660, 26057, 26054, 25242, 23980, 23175, 22757, 22701, 
    22922, 23356, 24334, 25235, 26457, 25509, 26713, 26682, 26112, 25469, 
    24752, 24205,
  24928, 24787, 26526, 26594, 26198, 25274, 23946, 23127, 22698, 22693, 
    22922, 23363, 24366, 25359, 26563, 26688, 27360, 26732, 26119, 25500, 
    24785, 24199,
  25636, 25513, 27104, 26876, 26326, 25293, 23914, 23166, 22719, 22765, 
    22971, 23483, 24152, 25513, 26556, 27298, 27479, 26813, 26195, 25500, 
    24740, 24186,
  26011, 25951, 27148, 26979, 26370, 25271, 23925, 23181, 22710, 22742, 
    22979, 23481, 24204, 25268, 26432, 27423, 27510, 26813, 26181, 25575, 
    24779, 24253,
  26014, 26033, 27112, 26974, 26407, 25271, 23918, 23166, 22780, 22742, 
    22937, 23501, 24295, 25417, 26549, 27423, 27542, 26900, 26299, 25631, 
    24887, 24246,
  25702, 25780, 27044, 26847, 26284, 25218, 23925, 23175, 22734, 22760, 
    22968, 23273, 24263, 25632, 26810, 27392, 27529, 26914, 26271, 25656, 
    24926, 24253,
  25144, 25239, 26776, 26616, 26141, 25187, 23894, 23149, 22813, 22788, 
    22909, 23402, 24313, 25464, 26801, 27231, 27592, 26965, 26306, 25781, 
    24970, 24287,
  24359, 24445, 25976, 26112, 25984, 25086, 23891, 23125, 22784, 22757, 
    22912, 23410, 24172, 25567, 26301, 26506, 27299, 26900, 26382, 25819, 
    25073, 24528,
  23334, 23426, 24896, 25455, 25651, 24999, 23794, 23134, 22822, 22795, 
    22869, 23420, 24153, 25495, 26806, 25416, 26476, 26770, 26389, 25949, 
    25009, 24502,
  22132, 22263, 23979, 24911, 25454, 24929, 23804, 23108, 22746, 22726, 
    22955, 23438, 24316, 25413, 26620, 24369, 25773, 26676, 26354, 25844, 
    25181, 24555,
  20950, 21124, 22996, 24389, 25205, 24817, 23776, 23079, 22747, 22755, 
    22955, 23447, 24136, 25353, 26387, 23154, 25113, 26619, 26321, 25863, 
    25124, 24569,
  20031, 20213, 22377, 23985, 25077, 24787, 23693, 23100, 22720, 22795, 
    22913, 23414, 24274, 25558, 26726, 22226, 24957, 26518, 26321, 25844, 
    25137, 24543,
  19482, 19648, 22355, 24018, 25057, 24820, 23725, 23070, 22759, 22750, 
    23009, 23419, 24304, 25486, 26528, 22078, 24696, 26547, 26293, 25894, 
    25175, 24637,
  19199, 19365, 23080, 24424, 25214, 24809, 23722, 23059, 22791, 22810, 
    23004, 23422, 24314, 25474, 26646, 23008, 25176, 26597, 26382, 25894, 
    25252, 24670,
  19000, 19185, 24136, 25030, 25398, 24829, 23684, 23085, 22797, 22767, 
    22925, 23427, 24314, 25598, 26594, 24395, 26576, 26706, 26328, 25888, 
    25252, 24617,
  18816, 18996, 24167, 25001, 25404, 24832, 23631, 23045, 22777, 22745, 
    22956, 23463, 24272, 25463, 26657, 24514, 26714, 26756, 26342, 25801, 
    25252, 24658,
  18729, 18854, 23103, 24486, 25198, 24743, 23645, 23021, 22748, 22774, 
    22996, 23412, 24344, 25510, 26487, 23051, 25500, 26634, 26328, 25845, 
    25145, 24645,
  18817, 18872, 22749, 24288, 25118, 24661, 23611, 23074, 22801, 22863, 
    23127, 23471, 24377, 25612, 26853, 22346, 25102, 26547, 26218, 25826, 
    25120, 24544,
  19001, 19029, 23251, 24514, 25226, 24678, 23604, 23037, 22854, 22843, 
    23019, 23522, 24441, 25451, 26976, 23259, 25893, 26613, 26232, 25751, 
    25152, 24652,
  19084, 19149, 23299, 24605, 25187, 24676, 23535, 23016, 22825, 22852, 
    23057, 23550, 24397, 25487, 26795, 23509, 25725, 26613, 26163, 25734, 
    25222, 24625,
  18953, 19086, 22937, 24377, 25106, 24575, 23529, 22996, 22790, 22809, 
    23006, 23568, 24368, 25575, 26814, 22737, 25295, 26476, 26198, 25697, 
    25120, 24625,
  18723, 18908, 22626, 24248, 25018, 24514, 23515, 22996, 22802, 22869, 
    22995, 23560, 24432, 25496, 26597, 22109, 25352, 26476, 26184, 25790, 
    25140, 24666,
  18654, 18847, 22692, 24289, 25021, 24531, 23487, 22979, 22817, 22878, 
    23012, 23462, 24575, 25529, 26507, 21856, 25451, 26432, 26129, 25728, 
    25064, 24512,
  18930, 19081, 22991, 24437, 25018, 24469, 23446, 22991, 22817, 22847, 
    23080, 23602, 24545, 25782, 27025, 22003, 25532, 26397, 26088, 25642, 
    24930, 24499,
  19524, 19594, 23589, 24695, 25116, 24383, 23422, 22970, 22799, 22911, 
    23092, 23505, 24514, 25772, 26647, 22462, 25669, 26376, 25999, 25505, 
    24898, 24392,
  20284, 20256, 24278, 25013, 25145, 24436, 23401, 22950, 22844, 22931, 
    23041, 23556, 24576, 25767, 26810, 23167, 25931, 26376, 25929, 25468, 
    24886, 24359,
  21095, 20986, 24651, 25228, 25211, 24383, 23388, 22953, 22818, 22905, 
    23093, 23635, 24553, 25837, 27029, 23741, 26118, 26360, 25978, 25499, 
    24893, 24427,
  21917, 21778, 24876, 25299, 25196, 24310, 23349, 22947, 22870, 22911, 
    23110, 23633, 24559, 25772, 26810, 23938, 26118, 26382, 25957, 25568, 
    24931, 24407,
  22649, 22557, 25089, 25401, 25151, 24294, 23329, 22972, 22839, 22923, 
    23042, 23646, 24643, 25804, 26839, 23848, 25913, 26398, 26026, 25637, 
    25002, 24508,
  23068, 23074, 25279, 25511, 25162, 24249, 23312, 22936, 22842, 22909, 
    23176, 23555, 24535, 25912, 27188, 23884, 25869, 26398, 26013, 25606, 
    25110, 24521,
  22956, 23060, 25348, 25549, 25148, 24210, 23225, 22919, 22822, 22921, 
    23108, 23725, 24644, 25979, 26639, 24235, 26056, 26312, 25938, 25525, 
    24926, 24481,
  22313, 22467, 25305, 25520, 25057, 24109, 23180, 22881, 22842, 22976, 
    23040, 23807, 24705, 26106, 26932, 24469, 26329, 26348, 25945, 25401, 
    24907, 24314,
  21405, 21498, 25006, 25399, 25008, 24037, 23195, 22902, 22831, 22956, 
    23154, 23809, 24868, 26217, 27060, 23760, 26250, 26348, 25959, 25526, 
    24952, 24382,
  20577, 20458, 24794, 25291, 24957, 24012, 23146, 22908, 22863, 22959, 
    23175, 23766, 24932, 26003, 27009, 22813, 26156, 26348, 25973, 25470, 
    24901, 24395,
  20051, 19650, 24953, 25278, 24886, 23937, 23115, 22846, 22826, 22922, 
    23217, 23713, 24871, 26207, 27162, 23073, 26101, 26298, 25898, 25433, 
    24838, 24275,
  19879, 19342, 25224, 25367, 24863, 23833, 23105, 22823, 22817, 22991, 
    23289, 23818, 24797, 26129, 27118, 23357, 26101, 26132, 25718, 25247, 
    24584, 24028,
  28696, 28660, 27792, 27110, 25741, 24124, 22696, 22170, 22069, 22506, 
    22925, 23571, 24561, 25737, 26500, 28629, 28850, 27795, 27132, 26463, 
    25474, 24560,
  28656, 28626, 27868, 27159, 25888, 24258, 22786, 22241, 22066, 22520, 
    22919, 23619, 24588, 25832, 26348, 28593, 28894, 27816, 27146, 26407, 
    25390, 24306,
  28565, 28557, 27917, 27248, 26013, 24359, 22858, 22261, 22130, 22517, 
    22910, 23508, 24514, 25637, 26781, 28570, 28770, 27751, 27110, 26407, 
    25365, 24312,
  28474, 28504, 27882, 27221, 26076, 24445, 22903, 22299, 22109, 22514, 
    22904, 23510, 24600, 25723, 26481, 28501, 28682, 27578, 27007, 26345, 
    25358, 24359,
  28403, 28474, 27838, 27213, 26122, 24515, 23007, 22304, 22106, 22456, 
    22929, 23570, 24489, 25835, 26539, 28385, 28482, 27499, 26882, 26232, 
    25345, 24412,
  28336, 28433, 27751, 27269, 26179, 24635, 23045, 22369, 22138, 22487, 
    22855, 23573, 24476, 25504, 26579, 28342, 28520, 27484, 26814, 26176, 
    25148, 24231,
  28267, 28364, 27726, 27276, 26256, 24691, 23114, 22386, 22143, 22407, 
    22812, 23469, 24316, 25478, 26449, 28347, 28471, 27542, 26814, 26065, 
    25001, 24010,
  28207, 28287, 27812, 27344, 26319, 24792, 23197, 22401, 22125, 22415, 
    22818, 23471, 24513, 25471, 26459, 28335, 28476, 27571, 26882, 26051, 
    25058, 24123,
  28161, 28230, 27843, 27406, 26341, 24833, 23249, 22521, 22169, 22449, 
    22826, 23364, 24350, 25710, 26429, 28347, 28551, 27585, 26785, 26001, 
    24988, 24016,
  28115, 28187, 27881, 27422, 26379, 24926, 23270, 22512, 22174, 22417, 
    22842, 23473, 24446, 25487, 26676, 28367, 28507, 27375, 26669, 25859, 
    24886, 24176,
  28047, 28121, 27739, 27379, 26460, 24962, 23336, 22550, 22192, 22454, 
    22822, 23384, 24458, 25729, 26504, 28260, 28332, 27173, 26496, 25846, 
    24924, 24135,
  27956, 28013, 27685, 27309, 26470, 24990, 23359, 22597, 22241, 22520, 
    22810, 23427, 24164, 25524, 26606, 28121, 28184, 27107, 26385, 25703, 
    24891, 24202,
  27870, 27893, 27604, 27244, 26429, 25037, 23446, 22579, 22282, 22448, 
    22759, 23439, 24221, 25449, 26550, 28007, 28053, 26841, 26144, 25535, 
    24732, 24195,
  27816, 27813, 27546, 27212, 26415, 25063, 23443, 22635, 22217, 22439, 
    22810, 23391, 24285, 25598, 26373, 27859, 27598, 26429, 25792, 25224, 
    24662, 23987,
  27792, 27783, 27376, 27126, 26341, 25009, 23522, 22664, 22267, 22464, 
    22792, 23310, 24082, 25314, 26687, 27692, 27187, 26141, 25667, 25187, 
    24502, 24081,
  27769, 27768, 27410, 27050, 26315, 25068, 23536, 22717, 22331, 22441, 
    22789, 23344, 24252, 25332, 26559, 27526, 27087, 26054, 25543, 25087, 
    24457, 24000,
  27722, 27722, 27343, 27072, 26372, 25163, 23591, 22734, 22304, 22473, 
    22821, 23337, 24244, 25402, 26679, 27296, 26894, 26054, 25619, 25099, 
    24476, 23886,
  27650, 27636, 27322, 27082, 26398, 25149, 23667, 22772, 22318, 22435, 
    22740, 23410, 24044, 25537, 26454, 27237, 26482, 26032, 25626, 25093, 
    24457, 23946,
  27566, 27534, 27360, 27187, 26446, 25235, 23681, 22793, 22342, 22449, 
    22766, 23361, 24125, 25295, 26588, 27396, 26906, 26054, 25660, 25055, 
    24463, 23879,
  27495, 27455, 27325, 27117, 26521, 25258, 23715, 22798, 22362, 22457, 
    22728, 23245, 24197, 25264, 26754, 27479, 26944, 25909, 25494, 24955, 
    24444, 23932,
  27466, 27421, 27322, 27117, 26535, 25339, 23754, 22875, 22403, 22503, 
    22791, 23303, 24093, 25422, 26573, 27479, 26987, 25895, 25459, 24980, 
    24450, 23865,
  27475, 27419, 27479, 27222, 26566, 25350, 23771, 22901, 22420, 22454, 
    22754, 23401, 24090, 25224, 26345, 27631, 27049, 26032, 25576, 25141, 
    24481, 23924,
  27470, 27408, 27447, 27187, 26529, 25333, 23764, 22924, 22393, 22474, 
    22830, 23399, 24236, 25399, 26420, 27759, 27104, 26067, 25507, 25073, 
    24443, 23938,
  27411, 27363, 27299, 27101, 26476, 25268, 23791, 22912, 22411, 22491, 
    22790, 23452, 24166, 25219, 26707, 27581, 27029, 26016, 25507, 25004, 
    24449, 23770,
  27332, 27305, 27188, 26960, 26400, 25302, 23868, 22933, 22416, 22482, 
    22790, 23276, 24257, 25296, 26568, 27403, 26893, 25944, 25493, 24942, 
    24366, 23864,
  27306, 27289, 27154, 27001, 26420, 25279, 23846, 22971, 22480, 22536, 
    22784, 23324, 24235, 25413, 26197, 27392, 26862, 25959, 25506, 24942, 
    24397, 23856,
  27356, 27343, 27337, 27039, 26425, 25301, 23895, 22956, 22498, 22504, 
    22773, 23322, 24069, 25438, 26129, 27509, 26868, 26051, 25596, 25010, 
    24448, 23937,
  27433, 27444, 27357, 27082, 26400, 25344, 23905, 22938, 22506, 22490, 
    22803, 23248, 24099, 25303, 26389, 27528, 26999, 26160, 25644, 25072, 
    24403, 23909,
  27473, 27518, 27299, 26957, 26365, 25315, 23891, 22965, 22483, 22490, 
    22721, 23334, 24064, 25375, 26529, 27434, 26954, 26196, 25699, 25158, 
    24409, 23949,
  27448, 27497, 27172, 26885, 26365, 25309, 23915, 23002, 22526, 22472, 
    22740, 23300, 24116, 25426, 26178, 27281, 26625, 26095, 25651, 25127, 
    24460, 23882,
  27345, 27355, 27104, 26847, 26296, 25250, 23922, 23023, 22503, 22521, 
    22829, 23308, 24199, 25065, 26526, 27150, 26463, 25950, 25512, 25096, 
    24511, 23889,
  27147, 27116, 27101, 26823, 26285, 25312, 23915, 23044, 22538, 22469, 
    22817, 23341, 24019, 25239, 26351, 26982, 26425, 25864, 25581, 25052, 
    24447, 24029,
  26853, 26818, 26923, 26774, 26304, 25317, 23974, 23076, 22541, 22495, 
    22794, 23328, 24192, 25311, 26347, 26921, 26088, 25763, 25471, 25039, 
    24453, 23988,
  26509, 26497, 26815, 26734, 26273, 25317, 23946, 23061, 22525, 22497, 
    22777, 23313, 24212, 25421, 26553, 26765, 25826, 25560, 25381, 24978, 
    24453, 24009,
  26199, 26198, 26617, 26610, 26204, 25343, 23977, 23075, 22569, 22534, 
    22820, 23356, 24288, 25379, 26487, 26587, 25701, 25430, 25236, 24958, 
    24414, 23968,
  25996, 25971, 26482, 26535, 26210, 25303, 23984, 23069, 22590, 22520, 
    22802, 23252, 24229, 25207, 26245, 26390, 25372, 25307, 25229, 24927, 
    24389, 23948,
  25922, 25853, 26441, 26529, 26179, 25320, 24005, 23108, 22616, 22537, 
    22853, 23376, 24196, 25439, 26154, 26217, 25198, 25170, 25077, 24883, 
    24471, 23907,
  25927, 25827, 26500, 26507, 26253, 25320, 23991, 23131, 22601, 22586, 
    22862, 23305, 24105, 25479, 26184, 26240, 25428, 25357, 25208, 24896, 
    24491, 23994,
  25917, 25809, 26624, 26529, 26250, 25345, 24053, 23125, 22601, 22571, 
    22825, 23226, 24127, 25376, 26295, 26376, 25832, 25545, 25422, 25051, 
    24503, 24095,
  25796, 25699, 26599, 26526, 26218, 25334, 24050, 23146, 22607, 22565, 
    22850, 23205, 24245, 25250, 26342, 26423, 25964, 25725, 25435, 25051, 
    24541, 24001,
  25526, 25445, 26507, 26432, 26173, 25362, 24057, 23151, 22583, 22562, 
    22816, 23355, 24004, 25297, 26363, 26254, 25814, 25639, 25373, 25020, 
    24503, 23987,
  25134, 25068, 26340, 26382, 26129, 25325, 24056, 23213, 22692, 22631, 
    22867, 23314, 24240, 25246, 26571, 26034, 25415, 25509, 25325, 24939, 
    24483, 24021,
  24715, 24651, 26001, 26165, 26084, 25300, 24018, 23157, 22645, 22606, 
    22822, 23256, 24183, 25192, 26079, 25735, 25048, 25328, 25297, 25026, 
    24611, 24081,
  24388, 24303, 25701, 26028, 26004, 25331, 24063, 23160, 22653, 22614, 
    22858, 23334, 24171, 25334, 26409, 25505, 24699, 25061, 25152, 24945, 
    24515, 24101,
  24235, 24107, 25642, 25995, 25946, 25322, 24032, 23181, 22689, 22602, 
    22841, 23388, 24062, 25421, 26266, 25480, 24904, 25198, 25214, 25013, 
    24643, 24027,
  24260, 24084, 25823, 26063, 26001, 25295, 24067, 23204, 22691, 22640, 
    22793, 23286, 24134, 25351, 26304, 25532, 25054, 25213, 25228, 24983, 
    24579, 24094,
  24399, 24200, 25764, 26041, 26026, 25300, 24067, 23175, 22683, 22568, 
    22827, 23375, 24178, 25378, 26157, 25452, 25041, 25328, 25304, 25044, 
    24604, 24155,
  24587, 24396, 25682, 26010, 26006, 25286, 24043, 23198, 22703, 22576, 
    22864, 23324, 24188, 25264, 26257, 25343, 25203, 25343, 25345, 25051, 
    24623, 24215,
  24775, 24604, 25762, 26051, 26018, 25306, 24043, 23166, 22712, 22582, 
    22804, 23373, 24218, 25381, 26465, 25502, 25701, 25595, 25462, 25181, 
    24604, 24155,
  24921, 24749, 25828, 26114, 26060, 25320, 24039, 23187, 22709, 22620, 
    22861, 23289, 24047, 25238, 26438, 25572, 25707, 25689, 25470, 25156, 
    24592, 24155,
  24970, 24773, 25875, 26106, 26047, 25337, 24029, 23151, 22686, 22631, 
    22819, 23395, 24146, 25320, 26514, 25663, 25615, 25523, 25393, 25094, 
    24573, 24208,
  24852, 24637, 25960, 26210, 26118, 25261, 24049, 23201, 22723, 22640, 
    22841, 23304, 24144, 25260, 26344, 25754, 25782, 25516, 25393, 25100, 
    24655, 24155,
  24519, 24316, 25909, 26151, 26078, 25289, 24008, 23166, 22715, 22674, 
    22796, 23236, 24149, 25157, 26441, 25682, 26013, 25646, 25435, 25100, 
    24604, 24121,
  23983, 23819, 25546, 25925, 25970, 25258, 24005, 23178, 22756, 22660, 
    22893, 23294, 24119, 25351, 26041, 25441, 26219, 25885, 25518, 25126, 
    24560, 24162,
  23338, 23220, 25072, 25650, 25843, 25261, 24036, 23184, 22738, 22651, 
    22827, 23433, 24171, 25390, 26646, 24953, 26444, 26129, 25663, 25181, 
    24687, 24108,
  22723, 22647, 24514, 25365, 25734, 25202, 24039, 23213, 22709, 22706, 
    22921, 23317, 24262, 25369, 26547, 24288, 26269, 26274, 25753, 25194, 
    24630, 24115,
  22258, 22205, 24456, 25300, 25709, 25200, 24008, 23178, 22738, 22651, 
    22888, 23310, 24243, 25279, 26468, 24001, 26095, 26325, 25774, 25219, 
    24554, 24115,
  22006, 21951, 24400, 25276, 25674, 25194, 24033, 23181, 22785, 22712, 
    22813, 23281, 24139, 25577, 26519, 24054, 26356, 26454, 25904, 25344, 
    24694, 24149,
  21994, 21912, 24481, 25322, 25709, 25155, 23963, 23196, 22759, 22726, 
    22899, 23279, 24142, 25414, 26698, 24157, 26200, 26535, 26022, 25362, 
    24726, 24149,
  22229, 22108, 24676, 25417, 25795, 25194, 23984, 23208, 22745, 22675, 
    22927, 23373, 24201, 25458, 26567, 24382, 26338, 26542, 26044, 25332, 
    24669, 24115,
  22676, 22519, 24963, 25637, 25864, 25203, 23963, 23179, 22730, 22640, 
    22959, 23414, 24226, 25320, 26526, 24853, 26375, 26629, 26037, 25363, 
    24720, 24202,
  23219, 23055, 25592, 25996, 25967, 25200, 23946, 23164, 22821, 22744, 
    22925, 23404, 24145, 25388, 26553, 25757, 26893, 26694, 26092, 25456, 
    24765, 24135,
  23691, 23563, 26154, 26362, 26126, 25214, 23946, 23152, 22754, 22732, 
    22919, 23338, 24365, 25489, 26410, 26590, 27404, 26831, 26244, 25518, 
    24873, 24250,
  23945, 23893, 26419, 26462, 26126, 25222, 23891, 23158, 22742, 22681, 
    22886, 23376, 24320, 25255, 26272, 26846, 27472, 26875, 26334, 25606, 
    24880, 24351,
  23929, 23970, 26323, 26429, 26122, 25163, 23933, 23158, 22719, 22721, 
    22977, 23412, 24175, 25358, 26119, 26857, 27516, 26962, 26320, 25704, 
    24931, 24351,
  23677, 23802, 25945, 26219, 26010, 25133, 23852, 23161, 22760, 22733, 
    22948, 23394, 24094, 25566, 26623, 26617, 27528, 26982, 26362, 25754, 
    25020, 24451,
  23242, 23420, 25389, 25851, 25821, 25108, 23874, 23162, 22778, 22736, 
    23014, 23407, 24333, 25228, 26354, 26029, 27254, 26853, 26376, 25785, 
    25084, 24378,
  22634, 22828, 24535, 25301, 25532, 24973, 23846, 23130, 22764, 22782, 
    22883, 23380, 24230, 25606, 26610, 24834, 26338, 26695, 26328, 25824, 
    25091, 24432,
  21824, 22019, 23813, 24787, 25361, 24909, 23843, 23112, 22781, 22774, 
    22952, 23293, 24304, 25575, 26321, 23698, 25360, 26579, 26341, 25837, 
    25104, 24398,
  20836, 21035, 23375, 24526, 25232, 24853, 23787, 23156, 22831, 22777, 
    22986, 23451, 24129, 25522, 26459, 23040, 25286, 26587, 26397, 25929, 
    25168, 24553,
  19819, 20014, 22792, 24203, 25135, 24803, 23773, 23101, 22802, 22769, 
    22984, 23509, 24311, 25427, 26579, 22425, 25074, 26535, 26382, 25904, 
    25302, 24573,
  18992, 19157, 22328, 23951, 25055, 24794, 23787, 23113, 22811, 22829, 
    22884, 23467, 24225, 25534, 26485, 21856, 24732, 26515, 26335, 25868, 
    25206, 24540,
  18485, 18617, 22169, 23821, 25020, 24781, 23718, 23086, 22820, 22812, 
    22984, 23396, 24319, 25555, 26628, 21680, 24726, 26529, 26404, 25881, 
    25226, 24614,
  18247, 18380, 22323, 23983, 25052, 24719, 23698, 23092, 22774, 22869, 
    22947, 23507, 24393, 25436, 26740, 22108, 24894, 26544, 26384, 25900, 
    25290, 24694,
  18115, 18288, 22777, 24285, 25121, 24725, 23684, 23087, 22751, 22770, 
    22962, 23467, 24248, 25522, 26557, 22952, 25417, 26573, 26329, 25900, 
    25220, 24635,
  17980, 18176, 22816, 24282, 25118, 24714, 23657, 23096, 22812, 22784, 
    22897, 23437, 24344, 25529, 26829, 22965, 25542, 26551, 26322, 25826, 
    25258, 24554,
  17849, 18015, 22380, 24040, 24993, 24621, 23605, 23026, 22797, 22781, 
    22957, 23483, 24298, 25565, 26595, 22163, 25138, 26544, 26176, 25782, 
    25208, 24695,
  17778, 17886, 22236, 24000, 24984, 24652, 23598, 23040, 22748, 22828, 
    23005, 23455, 24362, 25320, 26423, 21747, 25082, 26516, 26212, 25795, 
    25265, 24722,
  17759, 17836, 22327, 24035, 25007, 24627, 23588, 23041, 22822, 22868, 
    23057, 23435, 24353, 25800, 26748, 22048, 25219, 26501, 26267, 25839, 
    25138, 24749,
  17727, 17825, 22480, 24121, 25004, 24580, 23543, 23002, 22813, 22871, 
    23065, 23537, 24368, 25728, 26895, 22097, 25201, 26473, 26198, 25701, 
    25081, 24562,
  17675, 17823, 22477, 24084, 25005, 24541, 23504, 23038, 22772, 22831, 
    23068, 23542, 24314, 25598, 26610, 21846, 25263, 26473, 26123, 25671, 
    25100, 24596,
  17737, 17922, 22530, 24149, 25002, 24485, 23487, 23047, 22822, 22866, 
    23060, 23580, 24361, 25595, 26760, 21714, 25375, 26494, 26247, 25671, 
    25088, 24576,
  18099, 18274, 22749, 24286, 25033, 24471, 23470, 23009, 22811, 22858, 
    23066, 23558, 24412, 25882, 26922, 21805, 25494, 26479, 26165, 25653, 
    25031, 24583,
  18818, 18931, 23314, 24542, 25079, 24429, 23443, 23018, 22872, 22970, 
    23098, 23627, 24499, 25596, 27046, 22181, 25494, 26394, 26047, 25591, 
    24910, 24396,
  19754, 19773, 24097, 24878, 25165, 24471, 23454, 22975, 22867, 22938, 
    22998, 23592, 24440, 25845, 26637, 23003, 25835, 26300, 26006, 25548, 
    24802, 24262,
  20696, 20622, 24649, 25177, 25197, 24388, 23388, 22963, 22870, 22910, 
    23155, 23592, 24487, 25822, 26801, 23808, 26141, 26300, 25993, 25399, 
    24694, 24256,
  21541, 21408, 24895, 25304, 25180, 24352, 23395, 22948, 22859, 22956, 
    23195, 23572, 24544, 25754, 27123, 24167, 26228, 26344, 25931, 25486, 
    24879, 24350,
  22304, 22173, 24944, 25355, 25185, 24296, 23336, 22961, 22827, 22914, 
    23082, 23615, 24446, 25850, 26876, 24002, 26148, 26431, 25985, 25555, 
    25001, 24457,
  22961, 22893, 25045, 25369, 25120, 24268, 23284, 22902, 22833, 22960, 
    23182, 23659, 24594, 25659, 26938, 23762, 25943, 26366, 26028, 25598, 
    25033, 24551,
  23343, 23366, 25228, 25444, 25129, 24209, 23288, 22932, 22851, 22928, 
    23134, 23616, 24619, 26039, 26651, 23801, 25775, 26431, 26082, 25592, 
    25084, 24592,
  23254, 23355, 25382, 25504, 25078, 24148, 23254, 22897, 22798, 22963, 
    23120, 23687, 24695, 26026, 26831, 24305, 26110, 26401, 25979, 25587, 
    24913, 24331,
  22679, 22812, 25446, 25550, 25083, 24128, 23205, 22900, 22848, 23027, 
    23194, 23728, 24804, 25910, 26749, 24573, 26373, 26381, 25946, 25450, 
    24849, 24358,
  21826, 21900, 25106, 25377, 25021, 24103, 23185, 22921, 22837, 22987, 
    23206, 23746, 24762, 26121, 26940, 23978, 26354, 26331, 25987, 25500, 
    24868, 24419,
  20982, 20869, 24788, 25273, 24966, 24006, 23160, 22903, 22840, 22984, 
    23243, 23839, 24901, 26126, 27267, 22984, 26185, 26317, 25960, 25370, 
    24881, 24419,
  20382, 20023, 24899, 25243, 24861, 23924, 23088, 22895, 22858, 22973, 
    23183, 23771, 24837, 26014, 26800, 23062, 26249, 26273, 25932, 25451, 
    24926, 24386,
  20166, 19689, 25135, 25284, 24807, 23838, 23071, 22865, 22844, 22970, 
    23235, 23873, 24968, 26212, 27212, 23351, 26193, 26245, 25768, 25302, 
    24717, 24252,
  28681, 28618, 27874, 27042, 25766, 24118, 22715, 22191, 22080, 22506, 
    22866, 23602, 24691, 25874, 26272, 28669, 28881, 27825, 27201, 26439, 
    25568, 24540,
  28643, 28597, 27838, 27139, 25903, 24222, 22788, 22187, 22071, 22497, 
    22780, 23526, 24354, 25723, 26724, 28579, 28862, 27862, 27284, 26501, 
    25511, 24486,
  28561, 28555, 27919, 27220, 25994, 24373, 22857, 22270, 22155, 22499, 
    22922, 23584, 24474, 25795, 26554, 28585, 28893, 27869, 27166, 26476, 
    25479, 24526,
  28484, 28525, 27944, 27241, 26063, 24451, 22916, 22346, 22132, 22479, 
    22857, 23582, 24550, 25756, 26799, 28569, 28737, 27753, 27166, 26376, 
    25497, 24525,
  28423, 28499, 27838, 27235, 26143, 24526, 23019, 22345, 22128, 22536, 
    22902, 23482, 24432, 25679, 26842, 28440, 28551, 27515, 26882, 26190, 
    25242, 24304,
  28361, 28446, 27898, 27298, 26179, 24599, 23092, 22357, 22154, 22504, 
    22899, 23518, 24572, 25637, 26624, 28401, 28532, 27501, 26785, 26128, 
    25172, 24150,
  28285, 28353, 27807, 27290, 26297, 24714, 23158, 22430, 22186, 22504, 
    22770, 23464, 24480, 25673, 26641, 28314, 28538, 27565, 26882, 26157, 
    25108, 24150,
  28202, 28245, 27790, 27362, 26340, 24775, 23196, 22480, 22177, 22449, 
    22819, 23547, 24404, 25781, 26559, 28376, 28507, 27607, 26917, 26059, 
    25083, 24236,
  28121, 28152, 27812, 27332, 26360, 24873, 23265, 22494, 22209, 22460, 
    22838, 23542, 24520, 25676, 26549, 28312, 28476, 27572, 26814, 26082, 
    25038, 24176,
  28039, 28078, 27769, 27346, 26368, 24934, 23334, 22579, 22206, 22538, 
    22937, 23557, 24389, 25618, 26774, 28262, 28339, 27392, 26682, 25996, 
    24948, 24128,
  27945, 27992, 27701, 27292, 26385, 24957, 23376, 22576, 22197, 22468, 
    22732, 23468, 24319, 25499, 26751, 28120, 28114, 27103, 26462, 25816, 
    25031, 24363,
  27844, 27875, 27597, 27217, 26431, 24987, 23417, 22588, 22208, 22508, 
    22783, 23414, 24257, 25538, 26462, 27974, 27884, 26879, 26129, 25549, 
    24871, 24215,
  27764, 27758, 27528, 27126, 26391, 25066, 23455, 22620, 22234, 22405, 
    22772, 23452, 24173, 25468, 26796, 27851, 27710, 26540, 25909, 25343, 
    24692, 24074,
  27723, 27692, 27410, 27054, 26328, 25026, 23472, 22632, 22231, 22487, 
    22811, 23313, 24326, 25528, 26572, 27656, 27323, 26229, 25737, 25163, 
    24559, 24027,
  27708, 27682, 27274, 26969, 26304, 25037, 23514, 22663, 22260, 22473, 
    22820, 23307, 24301, 25577, 26476, 27394, 26937, 26028, 25571, 25162, 
    24552, 23866,
  27683, 27673, 27229, 26966, 26282, 25060, 23548, 22722, 22336, 22458, 
    22793, 23335, 24227, 25505, 26749, 27143, 26494, 25840, 25460, 25032, 
    24431, 23899,
  27622, 27608, 27259, 26976, 26299, 25084, 23614, 22766, 22367, 22467, 
    22836, 23405, 24246, 25351, 26454, 27143, 26550, 25912, 25557, 25050, 
    24557, 24079,
  27526, 27485, 27312, 27074, 26432, 25185, 23617, 22789, 22382, 22466, 
    22864, 23359, 24241, 25390, 26916, 27326, 26949, 26200, 25715, 25224, 
    24570, 23938,
  27422, 27351, 27235, 27103, 26435, 25244, 23683, 22807, 22358, 22460, 
    22844, 23324, 24177, 25381, 26449, 27442, 27285, 26315, 25750, 25236, 
    24570, 23931,
  27347, 27259, 27026, 26882, 26387, 25246, 23676, 22801, 22352, 22514, 
    22878, 23326, 24132, 25409, 26521, 27326, 27229, 26250, 25701, 25000, 
    24493, 23998,
  27329, 27230, 27129, 26954, 26419, 25283, 23745, 22874, 22372, 22500, 
    22795, 23321, 24270, 25371, 26410, 27360, 27142, 26099, 25542, 24987, 
    24410, 23897,
  27353, 27247, 27398, 27100, 26519, 25286, 23794, 22921, 22422, 22499, 
    22823, 23343, 24144, 25490, 26254, 27615, 27035, 25968, 25514, 24949, 
    24435, 23944,
  27367, 27267, 27347, 27089, 26490, 25319, 23801, 22900, 22424, 22459, 
    22780, 23303, 24282, 25513, 26582, 27682, 26860, 25788, 25335, 24868, 
    24352, 23890,
  27346, 27266, 27204, 27003, 26453, 25328, 23825, 22959, 22436, 22482, 
    22786, 23365, 24211, 25418, 26521, 27540, 26868, 25874, 25397, 24930, 
    24332, 23970,
  27321, 27262, 27179, 26954, 26450, 25341, 23880, 22929, 22486, 22461, 
    22802, 23277, 24163, 25443, 26322, 27456, 26979, 26047, 25589, 25104, 
    24498, 23809,
  27343, 27295, 27284, 27051, 26412, 25307, 23880, 22991, 22468, 22470, 
    22768, 23381, 24089, 25418, 26562, 27504, 27092, 26213, 25720, 25123, 
    24549, 23876,
  27410, 27380, 27292, 27085, 26467, 25336, 23904, 22988, 22497, 22467, 
    22905, 23337, 24032, 25492, 26462, 27548, 27079, 26256, 25762, 25153, 
    24447, 23956,
  27471, 27480, 27301, 26968, 26329, 25299, 23886, 22988, 22531, 22515, 
    22810, 23410, 24237, 25401, 26573, 27462, 26910, 26170, 25726, 25159, 
    24504, 23902,
  27486, 27531, 27210, 26903, 26338, 25254, 23879, 23014, 22549, 22486, 
    22850, 23408, 24027, 25366, 26268, 27323, 26860, 26184, 25706, 25215, 
    24529, 24069,
  27442, 27483, 27170, 26932, 26346, 25287, 23896, 23052, 22534, 22483, 
    22807, 23255, 24263, 25326, 26675, 27212, 26717, 26147, 25706, 25190, 
    24548, 23955,
  27328, 27325, 27129, 26887, 26326, 25282, 23931, 23058, 22557, 22512, 
    22847, 23298, 24189, 25342, 26493, 27156, 26704, 26132, 25720, 25122, 
    24535, 23961,
  27108, 27069, 27029, 26857, 26292, 25296, 23945, 23093, 22499, 22443, 
    22793, 23364, 24113, 25338, 26079, 27192, 26710, 26154, 25706, 25208, 
    24592, 23961,
  26766, 26728, 26984, 26801, 26340, 25312, 23931, 23096, 22537, 22543, 
    22838, 23420, 24090, 25293, 26657, 27098, 26742, 26226, 25754, 25227, 
    24637, 24028,
  26343, 26327, 26854, 26749, 26289, 25295, 23993, 23069, 22545, 22431, 
    22741, 23427, 24162, 25403, 26663, 27010, 26673, 26125, 25726, 25177, 
    24547, 24055,
  25938, 25926, 26657, 26614, 26235, 25326, 23993, 23087, 22592, 22563, 
    22824, 23252, 24117, 25307, 26375, 26857, 26374, 25901, 25595, 25164, 
    24591, 24115,
  25647, 25610, 26376, 26442, 26197, 25337, 24014, 23113, 22624, 22563, 
    22752, 23348, 24201, 25312, 26646, 26604, 26112, 25706, 25456, 25027, 
    24509, 24001,
  25519, 25443, 26246, 26428, 26182, 25337, 24011, 23131, 22621, 22543, 
    22857, 23229, 24223, 24990, 26110, 26451, 25963, 25562, 25353, 24953, 
    24540, 23980,
  25532, 25414, 26398, 26435, 26185, 25323, 23993, 23151, 22635, 22522, 
    22797, 23290, 24203, 25251, 26403, 26410, 25832, 25562, 25318, 24853, 
    24444, 24088,
  25591, 25438, 26431, 26576, 26203, 25376, 24069, 23181, 22632, 22508, 
    22849, 23305, 24147, 25300, 26071, 26532, 26087, 25676, 25353, 24978, 
    24514, 24067,
  25574, 25405, 26528, 26496, 26217, 25332, 24007, 23157, 22597, 22539, 
    22698, 23320, 24131, 25311, 26410, 26579, 26329, 25684, 25387, 24977, 
    24508, 23947,
  25399, 25242, 26365, 26447, 26151, 25329, 24021, 23136, 22664, 22548, 
    22794, 23236, 24138, 25223, 26672, 26435, 26218, 25691, 25346, 24896, 
    24438, 24000,
  25072, 24939, 26221, 26321, 26094, 25317, 24014, 23178, 22621, 22527, 
    22826, 23292, 24129, 25346, 26551, 26182, 25925, 25654, 25373, 24977, 
    24450, 24000,
  24681, 24556, 26057, 26221, 26068, 25233, 24045, 23157, 22697, 22587, 
    22829, 23320, 24250, 25283, 26296, 25901, 25588, 25475, 25324, 25002, 
    24489, 24047,
  24356, 24207, 25703, 26016, 25985, 25253, 24024, 23189, 22664, 22521, 
    22811, 23342, 24013, 25346, 26207, 25550, 25059, 25308, 25255, 24909, 
    24489, 24081,
  24188, 23999, 25515, 25929, 25957, 25295, 24038, 23207, 22714, 22567, 
    22771, 23162, 24173, 25328, 26401, 25391, 25077, 25250, 25200, 24996, 
    24565, 24141,
  24187, 23969, 25696, 25997, 26031, 25303, 24020, 23178, 22679, 22576, 
    22845, 23378, 24227, 25176, 26241, 25438, 25152, 25308, 25255, 25026, 
    24520, 24087,
  24302, 24080, 25769, 26046, 26016, 25317, 24031, 23192, 22725, 22613, 
    22865, 23355, 24264, 25160, 26560, 25502, 25239, 25395, 25339, 25014, 
    24501, 23973,
  24471, 24267, 25650, 26010, 26013, 25252, 24031, 23210, 22661, 22584, 
    22769, 23320, 24126, 25283, 26478, 25438, 25569, 25539, 25387, 24996, 
    24609, 24100,
  24649, 24464, 25647, 25981, 26004, 25236, 24044, 23189, 22699, 22639, 
    22886, 23286, 24126, 25388, 26267, 25491, 25676, 25539, 25408, 24983, 
    24539, 24047,
  24793, 24611, 25678, 26035, 26019, 25270, 24038, 23201, 22714, 22656, 
    22774, 23357, 24092, 25260, 26117, 25455, 25588, 25510, 25408, 25045, 
    24616, 24148,
  24850, 24657, 25751, 26046, 25999, 25298, 23992, 23198, 22679, 22596, 
    22851, 23271, 24128, 25325, 26362, 25519, 25731, 25597, 25435, 25045, 
    24565, 24208,
  24757, 24565, 25850, 26094, 26013, 25247, 24010, 23198, 22705, 22628, 
    22891, 23355, 24149, 25304, 26728, 25650, 25919, 25597, 25366, 24952, 
    24539, 24161,
  24466, 24304, 25782, 26089, 26051, 25295, 24003, 23181, 22728, 22622, 
    22811, 23368, 24126, 25395, 26132, 25653, 26193, 25792, 25477, 25033, 
    24571, 24107,
  23978, 23870, 25325, 25844, 25945, 25259, 23992, 23210, 22714, 22634, 
    22894, 23254, 24272, 25164, 26476, 25188, 26285, 25973, 25587, 25077, 
    24622, 24154,
  23366, 23316, 24679, 25448, 25750, 25216, 23979, 23151, 22755, 22628, 
    22937, 23353, 24223, 25521, 26343, 24372, 25950, 26110, 25601, 25107, 
    24559, 24000,
  22746, 22737, 24463, 25254, 25682, 25191, 23972, 23181, 22758, 22622, 
    22871, 23234, 24264, 25255, 26279, 23882, 25832, 26146, 25704, 25207, 
    24572, 24107,
  22201, 22201, 24567, 25359, 25726, 25197, 23989, 23216, 22711, 22645, 
    22857, 23279, 24050, 25246, 26389, 24115, 26237, 26356, 25863, 25288, 
    24622, 24134,
  21751, 21723, 24367, 25216, 25650, 25149, 23962, 23175, 22758, 22686, 
    22883, 23287, 24218, 25325, 26566, 24012, 26125, 26464, 25926, 25270, 
    24610, 24121,
  21388, 21312, 24147, 25117, 25642, 25107, 23975, 23178, 22743, 22711, 
    22812, 23338, 24122, 25377, 26491, 23772, 25856, 26479, 25960, 25345, 
    24661, 24162,
  21135, 21017, 24278, 25214, 25664, 25141, 23979, 23187, 22753, 22692, 
    22958, 23343, 24253, 25361, 26249, 24134, 26418, 26595, 26009, 25407, 
    24661, 24229,
  21041, 20900, 24200, 25133, 25604, 25130, 23923, 23184, 22741, 22668, 
    22880, 23277, 24186, 25302, 26676, 24226, 26274, 26660, 26092, 25519, 
    24770, 24188,
  21108, 20973, 24106, 25063, 25656, 25093, 23955, 23187, 22791, 22723, 
    22895, 23368, 24236, 25237, 26160, 24296, 26279, 26689, 26216, 25563, 
    24910, 24336,
  21258, 21161, 24195, 25128, 25607, 25138, 23931, 23187, 22800, 22632, 
    22904, 23313, 24339, 25358, 26823, 24599, 26299, 26703, 26237, 25650, 
    24885, 24316,
  21386, 21351, 24192, 25120, 25593, 25077, 23924, 23146, 22771, 22712, 
    22943, 23326, 24159, 25277, 26421, 24735, 26529, 26775, 26292, 25644, 
    24872, 24290,
  21428, 21473, 24038, 24983, 25525, 25035, 23882, 23199, 22812, 22712, 
    22929, 23379, 24142, 25316, 26343, 24526, 26162, 26775, 26389, 25725, 
    24962, 24384,
  21386, 21518, 23825, 24829, 25447, 25004, 23893, 23158, 22797, 22727, 
    22910, 23356, 24291, 25475, 26513, 24180, 25807, 26718, 26334, 25750, 
    24955, 24397,
  21279, 21476, 23661, 24694, 25353, 24962, 23855, 23120, 22768, 22770, 
    23001, 23334, 24254, 25499, 26493, 23851, 25321, 26668, 26403, 25868, 
    25052, 24425,
  21074, 21299, 23562, 24619, 25276, 24929, 23796, 23126, 22792, 22733, 
    22953, 23324, 24358, 25457, 26357, 23400, 25253, 26639, 26341, 25893, 
    25102, 24471,
  20696, 20921, 23446, 24593, 25288, 24887, 23800, 23135, 22769, 22807, 
    22999, 23378, 24273, 25587, 26797, 23102, 25241, 26545, 26341, 25881, 
    25269, 24505,
  20106, 20323, 23438, 24542, 25245, 24851, 23793, 23144, 22819, 22742, 
    22805, 23436, 24148, 25517, 26513, 23087, 25309, 26567, 26328, 25900, 
    25205, 24573,
  19381, 19583, 23146, 24383, 25188, 24828, 23768, 23150, 22781, 22757, 
    22945, 23416, 24383, 25184, 26821, 22770, 25216, 26524, 26354, 25782, 
    25167, 24660,
  18688, 18859, 22779, 24184, 25096, 24822, 23720, 23106, 22755, 22811, 
    22936, 23424, 24250, 25296, 26637, 22274, 25173, 26567, 26369, 25894, 
    25218, 24654,
  18163, 18300, 22371, 23979, 25071, 24761, 23689, 23095, 22755, 22746, 
    22857, 23416, 24262, 25676, 26196, 21869, 24942, 26538, 26314, 25875, 
    25250, 24627,
  17823, 17955, 22080, 23848, 24991, 24722, 23717, 23101, 22784, 22818, 
    22943, 23424, 24339, 25292, 26435, 21671, 24818, 26524, 26342, 25851, 
    25225, 24761,
  17580, 17744, 22005, 23819, 24939, 24711, 23689, 23107, 22790, 22800, 
    23000, 23483, 24317, 25320, 26390, 21707, 24775, 26495, 26232, 25770, 
    25295, 24661,
  17349, 17543, 22020, 23897, 24951, 24683, 23648, 23042, 22776, 22830, 
    22952, 23493, 24384, 25390, 26867, 21709, 24794, 26501, 26307, 25907, 
    25277, 24715,
  17120, 17303, 21962, 23800, 24959, 24658, 23631, 23116, 22838, 22816, 
    22926, 23488, 24350, 25404, 26395, 21502, 24862, 26590, 26239, 25807, 
    25207, 24668,
  16935, 17070, 22059, 23856, 24957, 24639, 23624, 23052, 22847, 22801, 
    23001, 23471, 24416, 25409, 26674, 21424, 25024, 26503, 26218, 25696, 
    25201, 24709,
  16824, 16915, 22145, 23911, 24940, 24602, 23593, 23070, 22806, 22810, 
    23001, 23529, 24340, 25511, 26737, 21512, 25168, 26446, 26156, 25696, 
    25169, 24649,
  16791, 16877, 22191, 24040, 24971, 24588, 23576, 23052, 22841, 22816, 
    23036, 23586, 24406, 25740, 26517, 21556, 25143, 26395, 26101, 25690, 
    25093, 24696,
  16892, 17011, 22320, 24073, 24980, 24530, 23521, 23053, 22827, 22854, 
    23138, 23550, 24353, 25665, 26846, 21625, 25286, 26482, 26116, 25709, 
    25239, 24683,
  17260, 17408, 22520, 24194, 24960, 24524, 23542, 23044, 22827, 22851, 
    23062, 23489, 24447, 25632, 26713, 21686, 25392, 26475, 26060, 25697, 
    25176, 24817,
  18009, 18139, 22832, 24347, 25035, 24511, 23500, 22956, 22854, 22834, 
    23048, 23536, 24459, 25647, 27217, 21939, 25337, 26381, 26006, 25585, 
    24947, 24469,
  19082, 19138, 23638, 24700, 25158, 24474, 23483, 23006, 22880, 22877, 
    23059, 23536, 24425, 25596, 26706, 22571, 25536, 26360, 26026, 25579, 
    24916, 24429,
  20240, 20204, 24457, 25061, 25166, 24444, 23434, 23003, 22846, 22926, 
    23022, 23531, 24566, 25835, 26624, 23530, 25897, 26345, 25972, 25431, 
    24878, 24369,
  21236, 21135, 24857, 25279, 25213, 24368, 23445, 23004, 22863, 22792, 
    23057, 23572, 24443, 25666, 26732, 24143, 26065, 26360, 25951, 25431, 
    24846, 24363,
  22001, 21884, 24868, 25308, 25213, 24343, 23393, 22978, 22869, 22927, 
    23137, 23587, 24505, 25925, 26745, 24178, 26090, 26274, 25951, 25469, 
    24885, 24443,
  22628, 22541, 24804, 25298, 25164, 24352, 23369, 22978, 22835, 22875, 
    23060, 23565, 24394, 25943, 26912, 23880, 26041, 26332, 25993, 25500, 
    24955, 24537,
  23174, 23141, 25002, 25414, 25159, 24305, 23366, 22955, 22850, 22908, 
    23172, 23643, 24552, 25697, 26532, 23826, 25892, 26339, 26035, 25525, 
    24968, 24611,
  23519, 23538, 25398, 25562, 25176, 24237, 23297, 22940, 22803, 22865, 
    23138, 23611, 24599, 26051, 26716, 24185, 25960, 26410, 26082, 25606, 
    25032, 24531,
  23475, 23532, 25547, 25565, 25107, 24145, 23224, 22902, 22844, 22931, 
    23144, 23697, 24749, 25909, 26876, 24612, 26147, 26404, 26035, 25531, 
    24988, 24445,
  22995, 23069, 25537, 25543, 25068, 24106, 23204, 22899, 22886, 22966, 
    23104, 23634, 24511, 26137, 26829, 24829, 26290, 26347, 25918, 25420, 
    24803, 24224,
  22221, 22248, 25271, 25374, 24999, 24011, 23207, 22864, 22848, 22958, 
    23147, 23678, 24686, 26072, 27046, 24257, 26316, 26275, 25953, 25377, 
    24835, 24398,
  21386, 21253, 24881, 25245, 24899, 23989, 23180, 22912, 22816, 22929, 
    23278, 23797, 24632, 26153, 26818, 23137, 26216, 26232, 25829, 25389, 
    24861, 24372,
  20735, 20384, 24874, 25216, 24836, 23908, 23083, 22865, 22825, 22921, 
    23188, 23810, 24790, 26032, 26929, 23003, 26104, 26189, 25760, 25315, 
    24747, 24198,
  20486, 20029, 25107, 25272, 24780, 23830, 23055, 22850, 22866, 22890, 
    23205, 23782, 24901, 26128, 27259, 23318, 26167, 26096, 25657, 25222, 
    24671, 24145,
  28647, 28573, 27862, 27073, 25763, 24167, 22678, 22216, 22137, 22487, 
    22920, 23628, 24608, 25588, 26746, 28588, 28810, 27896, 27197, 26440, 
    25499, 24460,
  28616, 28564, 27875, 27159, 25900, 24285, 22778, 22213, 22084, 22507, 
    22865, 23559, 24497, 25674, 26407, 28566, 28804, 27874, 27293, 26489, 
    25410, 24332,
  28547, 28548, 27929, 27185, 26014, 24383, 22843, 22281, 22122, 22435, 
    22851, 23576, 24659, 25792, 26431, 28563, 28842, 27860, 27182, 26432, 
    25410, 24372,
  28481, 28535, 27923, 27218, 26072, 24464, 22940, 22295, 22104, 22529, 
    22831, 23564, 24467, 25813, 26625, 28554, 28742, 27729, 27057, 26284, 
    25301, 24212,
  28427, 28507, 27887, 27323, 26140, 24595, 23013, 22357, 22136, 22480, 
    22899, 23500, 24472, 25725, 26545, 28454, 28512, 27571, 26824, 26122, 
    25060, 24098,
  28365, 28439, 27879, 27271, 26172, 24645, 23054, 22374, 22124, 22431, 
    22881, 23530, 24437, 25676, 26666, 28368, 28493, 27513, 26748, 25929, 
    24926, 24057,
  28281, 28322, 27807, 27263, 26279, 24754, 23124, 22421, 22170, 22474, 
    22872, 23391, 24385, 25601, 26607, 28340, 28443, 27549, 26810, 26010, 
    25002, 24063,
  28176, 28181, 27826, 27309, 26323, 24771, 23189, 22477, 22182, 22451, 
    22875, 23416, 24404, 25690, 26987, 28306, 28437, 27448, 26789, 26053, 
    24989, 24097,
  28057, 28045, 27747, 27282, 26351, 24852, 23227, 22494, 22190, 22474, 
    22743, 23438, 24422, 25689, 26295, 28242, 28318, 27224, 26554, 25910, 
    24969, 24103,
  27933, 27929, 27684, 27239, 26360, 24911, 23296, 22550, 22175, 22413, 
    22840, 23446, 24246, 25461, 26503, 28103, 28126, 27087, 26382, 25749, 
    24893, 24210,
  27811, 27817, 27570, 27198, 26334, 24944, 23365, 22531, 22222, 22501, 
    22860, 23359, 24275, 25496, 26556, 27969, 27870, 26784, 26132, 25475, 
    24886, 24189,
  27710, 27698, 27448, 27120, 26334, 24966, 23390, 22578, 22260, 22481, 
    22865, 23412, 24396, 25510, 26641, 27804, 27651, 26481, 25823, 25307, 
    24688, 24089,
  27653, 27600, 27351, 27047, 26279, 24974, 23414, 22601, 22201, 22467, 
    22862, 23432, 24238, 25575, 26728, 27570, 27322, 26213, 25643, 25121, 
    24453, 23941,
  27644, 27561, 27245, 26921, 26228, 24966, 23514, 22634, 22274, 22440, 
    22867, 23338, 24383, 25407, 26701, 27366, 26985, 26112, 25616, 25089, 
    24440, 23860,
  27648, 27572, 27147, 26879, 26168, 24977, 23521, 22675, 22332, 22466, 
    22790, 23434, 24280, 25632, 26897, 27012, 26332, 25903, 25471, 25020, 
    24370, 23894,
  27619, 27567, 27082, 26816, 26213, 25002, 23583, 22707, 22293, 22394, 
    22784, 23403, 24430, 25486, 26732, 26735, 25572, 25563, 25298, 24933, 
    24299, 23806,
  27536, 27489, 27081, 26899, 26229, 25083, 23604, 22760, 22334, 22491, 
    22827, 23342, 24202, 25383, 26795, 26885, 25801, 25628, 25401, 25001, 
    24439, 23940,
  27415, 27348, 27288, 26988, 26356, 25153, 23652, 22751, 22357, 22399, 
    22872, 23334, 24225, 25390, 26454, 27301, 26760, 26097, 25587, 25106, 
    24502, 23986,
  27295, 27206, 27132, 26969, 26388, 25212, 23663, 22803, 22345, 22379, 
    22937, 23435, 24365, 25534, 26451, 27378, 27184, 26291, 25697, 25131, 
    24534, 23953,
  27221, 27120, 26915, 26807, 26353, 25260, 23756, 22815, 22368, 22493, 
    22766, 23352, 24204, 25343, 26478, 27216, 27147, 26234, 25676, 25056, 
    24412, 23912,
  27213, 27101, 27070, 26917, 26388, 25217, 23742, 22900, 22386, 22421, 
    22797, 23356, 24172, 25474, 26698, 27344, 27203, 26190, 25607, 24969, 
    24355, 23825,
  27247, 27127, 27257, 27057, 26459, 25276, 23759, 22909, 22435, 22446, 
    22857, 23349, 24224, 25259, 26704, 27576, 27178, 26110, 25496, 25012, 
    24399, 23831,
  27277, 27164, 27226, 26974, 26459, 25270, 23780, 22912, 22423, 22475, 
    22686, 23277, 24221, 25368, 26223, 27610, 27091, 26125, 25530, 24950, 
    24316, 23784,
  27291, 27191, 27104, 26974, 26401, 25276, 23779, 22911, 22464, 22501, 
    22768, 23305, 24194, 25394, 26735, 27518, 27121, 26146, 25592, 24974, 
    24328, 23911,
  27318, 27218, 27176, 26998, 26404, 25267, 23831, 22961, 22458, 22409, 
    22834, 23328, 24181, 25350, 26610, 27515, 27078, 26218, 25606, 25111, 
    24481, 23850,
  27377, 27275, 27313, 27025, 26426, 25267, 23807, 22973, 22443, 22492, 
    22825, 23246, 24149, 25391, 26276, 27554, 27028, 26103, 25634, 25167, 
    24500, 23817,
  27441, 27368, 27254, 27057, 26418, 25325, 23873, 22964, 22513, 22497, 
    22876, 23325, 24195, 25372, 26584, 27513, 26947, 26081, 25599, 25092, 
    24398, 23917,
  27472, 27460, 27184, 26914, 26350, 25311, 23852, 22978, 22533, 22491, 
    22807, 23396, 24218, 25242, 26382, 27315, 26897, 26110, 25701, 25172, 
    24570, 23816,
  27454, 27492, 27169, 26901, 26324, 25297, 23886, 23037, 22516, 22525, 
    22858, 23365, 24249, 25282, 26194, 27282, 26791, 26203, 25729, 25172, 
    24480, 23970,
  27391, 27427, 27168, 26904, 26329, 25308, 23904, 23034, 22556, 22513, 
    22724, 23369, 24195, 25216, 26581, 27259, 26841, 26196, 25778, 25222, 
    24518, 23983,
  27262, 27257, 27100, 26887, 26285, 25297, 23914, 23016, 22524, 22476, 
    22713, 23286, 24126, 25274, 26560, 27248, 26784, 26116, 25653, 25141, 
    24524, 23916,
  27020, 26983, 27082, 26835, 26307, 25319, 23956, 23084, 22562, 22496, 
    22764, 23346, 24217, 25335, 26581, 27209, 26872, 26151, 25764, 25234, 
    24562, 24003,
  26638, 26605, 26963, 26766, 26272, 25272, 23938, 23101, 22568, 22527, 
    22769, 23314, 24347, 25277, 26448, 27206, 26859, 26231, 25729, 25171, 
    24569, 24049,
  26159, 26143, 26854, 26720, 26257, 25283, 23983, 23098, 22612, 22527, 
    22857, 23288, 24180, 25383, 26600, 27109, 26840, 26246, 25798, 25234, 
    24587, 24103,
  25683, 25672, 26659, 26612, 26192, 25300, 23976, 23148, 22570, 22544, 
    22789, 23278, 24157, 25358, 26464, 26967, 26747, 26101, 25687, 25090, 
    24517, 23968,
  25316, 25297, 26506, 26501, 26209, 25266, 23983, 23116, 22585, 22576, 
    22880, 23394, 24132, 25265, 26273, 26850, 26497, 25914, 25494, 25066, 
    24530, 23948,
  25129, 25089, 26321, 26410, 26129, 25291, 24021, 23148, 22617, 22595, 
    22848, 23404, 24034, 25509, 26624, 26669, 26174, 25653, 25335, 24903, 
    24377, 23988,
  25127, 25042, 26226, 26370, 26148, 25291, 24014, 23124, 22614, 22633, 
    22820, 23275, 24214, 25318, 26450, 26476, 25879, 25429, 25183, 24829, 
    24351, 23901,
  25230, 25080, 26184, 26324, 26114, 25310, 24000, 23156, 22614, 22616, 
    22868, 23374, 24229, 25376, 26268, 26399, 25918, 25444, 25155, 24785, 
    24364, 23914,
  25303, 25101, 26184, 26267, 26129, 25319, 24042, 23133, 22707, 22572, 
    22825, 23384, 24159, 25395, 26159, 26379, 25999, 25408, 25079, 24717, 
    24332, 23760,
  25229, 25025, 26174, 26285, 26128, 25310, 24024, 23165, 22663, 22575, 
    22811, 23320, 24071, 25353, 26244, 26338, 26185, 25552, 25238, 24804, 
    24434, 24008,
  24986, 24810, 26098, 26243, 26094, 25274, 24041, 23141, 22675, 22586, 
    22822, 23294, 24115, 25320, 26357, 26220, 26260, 25747, 25376, 24909, 
    24408, 24021,
  24654, 24492, 25945, 26135, 26014, 25257, 24031, 23174, 22634, 22583, 
    22879, 23333, 24198, 25267, 26544, 25984, 25768, 25601, 25320, 25040, 
    24484, 23994,
  24359, 24182, 25694, 25966, 25934, 25282, 24021, 23197, 22701, 22609, 
    22876, 23305, 24391, 25327, 26257, 25625, 25164, 25263, 25168, 24965, 
    24516, 24014,
  24196, 23995, 25491, 25896, 25904, 25243, 24055, 23171, 22707, 22595, 
    22828, 23363, 24157, 25238, 26478, 25377, 25114, 25154, 25099, 24809, 
    24433, 23974,
  24183, 23975, 25512, 25976, 25897, 25221, 24014, 23177, 22681, 22586, 
    22802, 23317, 24067, 25248, 26629, 25377, 25319, 25284, 25244, 24940, 
    24452, 24068,
  24279, 24082, 25732, 26009, 26014, 25288, 24014, 23168, 22666, 22534, 
    22868, 23350, 24206, 25294, 26689, 25477, 25612, 25371, 25259, 24990, 
    24446, 24101,
  24433, 24254, 25714, 26060, 26014, 25282, 24007, 23189, 22701, 22603, 
    22862, 23416, 24045, 25175, 26406, 25519, 25681, 25508, 25348, 24990, 
    24459, 24041,
  24600, 24435, 25684, 26017, 25988, 25254, 24058, 23162, 22669, 22661, 
    22888, 23305, 24018, 25227, 26488, 25457, 25662, 25494, 25320, 24978, 
    24580, 24081,
  24742, 24582, 25862, 26095, 25994, 25277, 24021, 23203, 22689, 22641, 
    22911, 23289, 24070, 25380, 26469, 25580, 25681, 25552, 25328, 25021, 
    24478, 24041,
  24810, 24656, 25915, 26170, 26014, 25310, 24045, 23203, 22716, 22692, 
    22913, 23350, 24169, 25278, 26501, 25660, 25998, 25601, 25369, 25083, 
    24522, 24061,
  24754, 24621, 25841, 26129, 26054, 25319, 24010, 23200, 22736, 22635, 
    22968, 23401, 24088, 25285, 26490, 25689, 26129, 25703, 25362, 24953, 
    24541, 24075,
  24536, 24444, 25748, 26095, 26022, 25268, 24014, 23159, 22721, 22712, 
    22990, 23383, 24208, 25444, 26285, 25644, 26329, 25862, 25466, 24959, 
    24497, 24021,
  24151, 24110, 25623, 26001, 26004, 25251, 23993, 23198, 22745, 22693, 
    22959, 23376, 24267, 25357, 26357, 25388, 26528, 26007, 25528, 25102, 
    24446, 24082,
  23635, 23645, 25162, 25753, 25876, 25266, 24007, 23198, 22733, 22727, 
    22976, 23389, 24174, 25388, 26551, 24770, 26217, 26166, 25673, 25102, 
    24586, 24155,
  23047, 23091, 24911, 25588, 25813, 25210, 23996, 23206, 22772, 22687, 
    22928, 23447, 24174, 25385, 26307, 24415, 26167, 26274, 25721, 25208, 
    24586, 24169,
  22413, 22459, 24900, 25570, 25825, 25201, 24017, 23218, 22772, 22756, 
    22817, 23376, 24214, 25390, 26410, 24561, 26503, 26412, 25832, 25239, 
    24638, 24175,
  21711, 21727, 24611, 25376, 25716, 25201, 24004, 23169, 22733, 22633, 
    23034, 23391, 24260, 25376, 26965, 24288, 26410, 26498, 25901, 25351, 
    24669, 24102,
  20928, 20905, 24203, 25128, 25642, 25165, 23972, 23189, 22769, 22721, 
    23005, 23379, 24236, 25253, 26435, 23858, 26085, 26535, 26004, 25345, 
    24676, 24156,
  20133, 20085, 23904, 24910, 25548, 25129, 23910, 23169, 22778, 22733, 
    22980, 23397, 24270, 25421, 26469, 23822, 26317, 26643, 26087, 25525, 
    24733, 24236,
  19471, 19415, 23243, 24549, 25384, 25061, 23920, 23163, 22763, 22708, 
    22974, 23343, 24209, 25586, 26278, 23257, 26124, 26622, 26204, 25538, 
    24925, 24297,
  19062, 19009, 22688, 24186, 25236, 25025, 23955, 23172, 22755, 22733, 
    22983, 23397, 24310, 25479, 26590, 22588, 25588, 26614, 26198, 25619, 
    24835, 24370,
  18923, 18881, 22363, 23995, 25121, 24983, 23879, 23172, 22731, 22728, 
    22906, 23293, 24148, 25482, 26484, 22349, 25220, 26615, 26232, 25688, 
    24919, 24243,
  18985, 18967, 22391, 23963, 25059, 24944, 23886, 23128, 22804, 22760, 
    22934, 23427, 24207, 25439, 26278, 22245, 24890, 26585, 26254, 25725, 
    24932, 24411,
  19170, 19199, 22381, 23936, 25027, 24876, 23869, 23172, 22767, 22751, 
    22980, 23435, 24170, 25193, 26535, 22192, 24729, 26449, 26281, 25707, 
    25002, 24431,
  19434, 19528, 22496, 23987, 25016, 24888, 23855, 23140, 22799, 22783, 
    22983, 23382, 24259, 25405, 26604, 22319, 24866, 26543, 26295, 25806, 
    25085, 24512,
  19740, 19893, 22800, 24184, 25133, 24888, 23817, 23120, 22761, 22772, 
    23058, 23337, 24432, 25337, 26423, 22542, 25090, 26579, 26406, 25875, 
    25117, 24633,
  20001, 20185, 23234, 24448, 25202, 24877, 23838, 23102, 22791, 22780, 
    23063, 23426, 24259, 25449, 26626, 22920, 25320, 26572, 26385, 25925, 
    25142, 24499,
  20091, 20285, 23571, 24620, 25288, 24866, 23779, 23117, 22738, 22749, 
    23009, 23540, 24289, 25573, 26416, 23257, 25532, 26615, 26379, 25981, 
    25244, 24633,
  19918, 20124, 23678, 24693, 25265, 24858, 23807, 23117, 22806, 22786, 
    23021, 23558, 24213, 25349, 26601, 23393, 25645, 26615, 26337, 25832, 
    25194, 24640,
  19499, 19723, 23510, 24620, 25216, 24774, 23751, 23094, 22771, 22764, 
    23004, 23462, 24400, 25482, 26649, 23195, 25570, 26522, 26331, 25807, 
    25188, 24493,
  18954, 19177, 23179, 24457, 25137, 24813, 23752, 23070, 22768, 22819, 
    23042, 23455, 24324, 25717, 26601, 22830, 25421, 26529, 26310, 25845, 
    25232, 24634,
  18415, 18610, 22680, 24161, 25062, 24760, 23728, 23115, 22800, 22781, 
    23028, 23475, 24366, 25564, 26426, 22267, 25240, 26522, 26282, 25913, 
    25284, 24694,
  17948, 18112, 22312, 23921, 24973, 24695, 23696, 23068, 22803, 22819, 
    22885, 23429, 24295, 25387, 26704, 21681, 24730, 26443, 26296, 25776, 
    25239, 24540,
  17540, 17701, 22102, 23830, 24942, 24693, 23700, 23091, 22810, 22810, 
    23065, 23597, 24384, 25603, 26831, 21433, 24593, 26457, 26200, 25801, 
    25157, 24534,
  17153, 17333, 21981, 23820, 24934, 24721, 23673, 23098, 22833, 22879, 
    23031, 23529, 24374, 25629, 26879, 21276, 24693, 26500, 26235, 25759, 
    25151, 24735,
  16788, 16973, 21918, 23784, 24911, 24626, 23634, 23071, 22848, 22865, 
    23180, 23585, 24360, 25488, 26501, 21290, 24843, 26465, 26151, 25715, 
    25087, 24668,
  16490, 16643, 21958, 23823, 24954, 24595, 23628, 23025, 22840, 22866, 
    23091, 23458, 24483, 25537, 26524, 21295, 24974, 26479, 26151, 25628, 
    25132, 24468,
  16312, 16412, 22106, 23849, 24957, 24587, 23593, 23063, 22823, 22838, 
    23103, 23497, 24439, 25718, 26807, 21366, 25074, 26435, 26098, 25685, 
    25107, 24569,
  16302, 16374, 22195, 23912, 24920, 24545, 23548, 23052, 22855, 22872, 
    23095, 23515, 24425, 25497, 26935, 21455, 25074, 26479, 26167, 25753, 
    25177, 24669,
  16545, 16634, 22311, 23998, 24963, 24542, 23538, 23005, 22846, 22835, 
    23052, 23578, 24514, 25772, 26996, 21569, 25273, 26479, 26174, 25760, 
    25209, 24689,
  17166, 17276, 22616, 24194, 24978, 24531, 23542, 23019, 22835, 22875, 
    23112, 23591, 24548, 25726, 26839, 21718, 25323, 26457, 26139, 25692, 
    25076, 24596,
  18212, 18293, 23125, 24464, 25072, 24520, 23507, 23041, 22891, 22899, 
    23030, 23632, 24541, 25951, 27195, 22111, 25379, 26387, 26050, 25592, 
    24974, 24476,
  19530, 19526, 23989, 24889, 25133, 24470, 23466, 23005, 22856, 22933, 
    23144, 23610, 24519, 25829, 27076, 23025, 25653, 26445, 26064, 25610, 
    24981, 24402,
  20802, 20712, 24699, 25217, 25210, 24456, 23463, 23000, 22886, 22939, 
    23170, 23595, 24591, 25754, 26897, 23900, 25990, 26416, 26057, 25629, 
    24968, 24490,
  21764, 21641, 24919, 25339, 25230, 24409, 23480, 22944, 22918, 22954, 
    23037, 23635, 24507, 25882, 26707, 24229, 25959, 26394, 26023, 25537, 
    24912, 24410,
  22393, 22296, 24762, 25255, 25167, 24333, 23421, 22989, 22883, 22943, 
    23213, 23575, 24544, 25978, 26822, 23958, 25940, 26344, 26001, 25469, 
    24937, 24417,
  22858, 22811, 24730, 25283, 25159, 24275, 23362, 22966, 22860, 22955, 
    23285, 23621, 24485, 26120, 27234, 23767, 25822, 26344, 25975, 25631, 
    25059, 24624,
  23288, 23275, 25158, 25522, 25176, 24255, 23366, 22945, 22837, 22926, 
    23180, 23773, 24621, 25910, 26992, 24258, 26257, 26359, 25941, 25600, 
    24995, 24471,
  23604, 23602, 25657, 25681, 25219, 24298, 23311, 22966, 22884, 23004, 
    23183, 23796, 24651, 25931, 27057, 24880, 26438, 26401, 26003, 25538, 
    24976, 24498,
  23620, 23629, 25695, 25681, 25168, 24141, 23290, 22951, 22829, 22967, 
    23109, 23718, 24676, 26022, 26882, 25204, 26432, 26345, 26003, 25600, 
    24913, 24338,
  23251, 23279, 25620, 25603, 25065, 24113, 23221, 22919, 22872, 22964, 
    23155, 23685, 24735, 26162, 27053, 25192, 26414, 26301, 25914, 25427, 
    24824, 24251,
  22577, 22578, 25315, 25439, 24980, 24060, 23170, 22914, 22879, 22930, 
    23215, 23794, 24790, 26197, 27031, 24589, 26420, 26237, 25832, 25377, 
    24761, 24218,
  21775, 21636, 24905, 25243, 24905, 23990, 23145, 22864, 22873, 22954, 
    23155, 23729, 24733, 26274, 26907, 23338, 26203, 26179, 25804, 25403, 
    24742, 24278,
  21099, 20756, 24865, 25200, 24825, 23929, 23111, 22885, 22859, 22968, 
    23264, 23830, 24832, 26307, 26770, 22999, 26110, 26129, 25729, 25366, 
    24711, 24232,
  20830, 20386, 25065, 25260, 24774, 23848, 23080, 22882, 22842, 22966, 
    23207, 23787, 24891, 26257, 27034, 23381, 26209, 26057, 25604, 25124, 
    24521, 23979,
  28614, 28535, 27829, 27110, 25779, 24131, 22728, 22194, 22107, 22516, 
    22849, 23655, 24587, 25679, 26781, 28625, 28940, 27901, 27285, 26544, 
    25417, 24433,
  28589, 28532, 27850, 27191, 25909, 24274, 22783, 22261, 22127, 22427, 
    22946, 23564, 24462, 25693, 26675, 28588, 28878, 27895, 27235, 26457, 
    25430, 24459,
  28534, 28525, 27857, 27215, 26003, 24341, 22849, 22272, 22121, 22455, 
    22940, 23531, 24609, 25801, 26829, 28579, 28791, 27801, 27167, 26457, 
    25353, 24332,
  28477, 28514, 27895, 27239, 26076, 24490, 22984, 22310, 22121, 22461, 
    22851, 23490, 24530, 25474, 26479, 28594, 28691, 27707, 27015, 26295, 
    25239, 24258,
  28421, 28481, 27850, 27279, 26132, 24553, 23012, 22328, 22118, 22472, 
    22811, 23568, 24409, 25743, 26679, 28496, 28548, 27635, 26946, 26165, 
    25035, 24245,
  28351, 28406, 27794, 27234, 26157, 24685, 23095, 22404, 22155, 22454, 
    22842, 23542, 24552, 25564, 26518, 28396, 28492, 27512, 26779, 26015, 
    24958, 24071,
  28251, 28279, 27735, 27325, 26209, 24702, 23129, 22416, 22161, 22445, 
    22845, 23413, 24386, 25666, 26515, 28343, 28367, 27432, 26656, 26015, 
    24945, 24084,
  28116, 28113, 27718, 27268, 26309, 24780, 23209, 22498, 22172, 22448, 
    22813, 23418, 24398, 25531, 26626, 28317, 28242, 27209, 26449, 25723, 
    24844, 23950,
  27955, 27934, 27654, 27254, 26309, 24830, 23264, 22503, 22178, 22433, 
    22822, 23400, 24300, 25489, 26670, 28206, 28143, 26942, 26270, 25629, 
    24716, 24043,
  27788, 27768, 27557, 27174, 26288, 24861, 23267, 22536, 22239, 22450, 
    22759, 23524, 24344, 25478, 26795, 28024, 27900, 26782, 26173, 25455, 
    24824, 24062,
  27646, 27628, 27357, 27013, 26246, 24869, 23333, 22565, 22259, 22502, 
    22741, 23483, 24169, 25617, 26640, 27756, 27514, 26423, 25849, 25343, 
    24626, 24055,
  27557, 27517, 27228, 26848, 26182, 24917, 23423, 22602, 22291, 22452, 
    22829, 23421, 24383, 25624, 26831, 27382, 27121, 26141, 25607, 25088, 
    24505, 23795,
  27538, 27454, 27142, 26810, 26148, 24874, 23436, 22644, 22241, 22412, 
    22815, 23396, 24400, 25381, 26347, 27145, 26269, 25824, 25407, 25001, 
    24397, 23888,
  27572, 27453, 27134, 26829, 26131, 24963, 23482, 22676, 22296, 22492, 
    22877, 23487, 24257, 25423, 26376, 27000, 26306, 25824, 25455, 25025, 
    24359, 23935,
  27602, 27487, 27076, 26789, 26188, 24966, 23481, 22720, 22346, 22429, 
    22831, 23451, 24427, 25498, 26582, 26891, 26007, 25779, 25483, 25007, 
    24422, 23887,
  27573, 27485, 27053, 26749, 26165, 25014, 23551, 22740, 22313, 22397, 
    22825, 23388, 24293, 25162, 26510, 26710, 25484, 25433, 25289, 24876, 
    24371, 23720,
  27475, 27400, 27124, 26818, 26245, 25098, 23603, 22716, 22351, 22448, 
    22828, 23420, 24187, 25616, 26229, 26828, 25484, 25368, 25282, 25006, 
    24440, 23967,
  27339, 27257, 27151, 26942, 26331, 25167, 23644, 22766, 22339, 22459, 
    22771, 23425, 24150, 25178, 26810, 27216, 26554, 25945, 25571, 25130, 
    24529, 23900,
  27215, 27126, 26967, 26867, 26299, 25145, 23675, 22757, 22377, 22477, 
    22787, 23354, 24157, 25232, 26472, 27263, 27214, 26241, 25757, 25055, 
    24535, 24033,
  27146, 27057, 26851, 26797, 26313, 25162, 23692, 22836, 22423, 22459, 
    22824, 23336, 24223, 25411, 26607, 27132, 27239, 26248, 25626, 25024, 
    24420, 23906,
  27139, 27052, 27053, 26872, 26342, 25190, 23744, 22907, 22449, 22496, 
    22816, 23368, 24223, 25360, 26346, 27364, 27146, 26118, 25550, 25055, 
    24363, 23838,
  27165, 27082, 27204, 26987, 26326, 25223, 23744, 22901, 22414, 22473, 
    22684, 23300, 24097, 25187, 26709, 27506, 26890, 25995, 25515, 25005, 
    24388, 23805,
  27191, 27121, 27159, 26901, 26353, 25228, 23796, 22871, 22437, 22461, 
    22789, 23409, 24333, 25306, 26695, 27531, 26684, 25894, 25474, 24948, 
    24381, 23844,
  27226, 27153, 27062, 26891, 26321, 25304, 23792, 22918, 22446, 22555, 
    22869, 23426, 24176, 25247, 26378, 27473, 26641, 25907, 25529, 25103, 
    24412, 23878,
  27292, 27187, 27149, 26934, 26350, 25250, 23796, 22938, 22469, 22423, 
    22806, 23317, 24202, 25445, 26167, 27523, 26815, 26074, 25618, 25141, 
    24489, 23897,
  27379, 27248, 27260, 27076, 26413, 25287, 23844, 22991, 22510, 22460, 
    22823, 23388, 24242, 25222, 26479, 27641, 27095, 26304, 25784, 25271, 
    24539, 23931,
  27444, 27339, 27232, 27032, 26404, 25287, 23868, 22982, 22469, 22472, 
    22774, 23304, 24121, 25268, 26394, 27560, 27157, 26319, 25825, 25165, 
    24545, 23944,
  27454, 27423, 27187, 26971, 26332, 25247, 23896, 23029, 22521, 22500, 
    22868, 23364, 24115, 25256, 26672, 27435, 26951, 26348, 25810, 25277, 
    24551, 23997,
  27412, 27442, 27151, 26917, 26307, 25262, 23878, 23032, 22518, 22546, 
    22728, 23258, 24115, 25329, 26656, 27376, 26901, 26247, 25845, 25283, 
    24570, 24097,
  27325, 27361, 27123, 26879, 26307, 25284, 23871, 23032, 22535, 22531, 
    22873, 23341, 24241, 25253, 26425, 27273, 26976, 26449, 25845, 25258, 
    24615, 24211,
  27169, 27173, 27123, 26863, 26298, 25250, 23912, 23058, 22550, 22540, 
    22899, 23257, 24162, 25440, 26707, 27262, 26901, 26332, 25893, 25357, 
    24653, 23989,
  26897, 26877, 27073, 26895, 26278, 25284, 23919, 23058, 22541, 22479, 
    22836, 23308, 24184, 25347, 26256, 27259, 26920, 26332, 25928, 25313, 
    24620, 24063,
  26490, 26470, 26978, 26807, 26269, 25272, 23951, 23081, 22614, 22536, 
    22822, 23277, 24075, 25153, 26679, 27181, 26865, 26325, 25954, 25319, 
    24633, 24116,
  25992, 25980, 26676, 26669, 26163, 25258, 23985, 23084, 22575, 22536, 
    22813, 23353, 24023, 25344, 26212, 27067, 26751, 26289, 25893, 25413, 
    24703, 24109,
  25495, 25491, 26567, 26535, 26126, 25255, 23978, 23057, 22584, 22550, 
    22870, 23259, 24352, 25318, 26476, 26997, 26726, 26304, 25920, 25406, 
    24684, 24210,
  25095, 25108, 26443, 26400, 26097, 25286, 23988, 23116, 22657, 22650, 
    22827, 23330, 24198, 25320, 26541, 26849, 26534, 26085, 25671, 25244, 
    24639, 24109,
  24869, 24893, 26226, 26373, 26049, 25246, 24020, 23116, 22654, 22532, 
    22775, 23292, 24134, 25313, 26415, 26671, 26185, 25625, 25416, 24996, 
    24531, 24022,
  24844, 24833, 26151, 26241, 26074, 25261, 23995, 23137, 22663, 22578, 
    22846, 23315, 24173, 25265, 26299, 26418, 25729, 25278, 25105, 24784, 
    24384, 23935,
  24961, 24866, 26042, 26222, 26063, 25277, 24006, 23142, 22668, 22650, 
    22844, 23317, 24161, 25306, 26426, 26201, 25487, 25176, 25009, 24753, 
    24269, 23868,
  25084, 24908, 26040, 26219, 26057, 25286, 24013, 23169, 22628, 22607, 
    22915, 23335, 24129, 25241, 26795, 26123, 25643, 25343, 25140, 24821, 
    24307, 23821,
  25081, 24880, 26062, 26238, 26114, 25328, 24006, 23204, 22680, 22621, 
    22798, 23355, 24104, 25195, 26282, 26131, 26035, 25667, 25416, 25014, 
    24479, 23981,
  24912, 24729, 25959, 26165, 26040, 25300, 23998, 23181, 22686, 22584, 
    22860, 23210, 24131, 25180, 26764, 26120, 26484, 25949, 25581, 25088, 
    24466, 23941,
  24642, 24475, 25819, 26101, 26106, 25308, 24037, 23186, 22753, 22658, 
    22889, 23350, 24166, 25481, 26139, 25956, 26409, 25899, 25478, 24989, 
    24543, 24008,
  24391, 24222, 25782, 26090, 26026, 25339, 24040, 23178, 22698, 22592, 
    22926, 23312, 24079, 25355, 26351, 25760, 26253, 25790, 25505, 25082, 
    24511, 24108,
  24248, 24077, 25621, 25987, 26031, 25272, 24050, 23183, 22689, 22595, 
    22823, 23261, 24148, 25229, 26265, 25538, 26141, 25768, 25457, 25076, 
    24562, 24061,
  24235, 24072, 25517, 25901, 25985, 25252, 24019, 23159, 22671, 22610, 
    22895, 23360, 24156, 25337, 26422, 25399, 26091, 25776, 25498, 25094, 
    24612, 24068,
  24318, 24168, 25606, 25944, 25974, 25316, 24047, 23204, 22715, 22649, 
    22854, 23317, 24094, 25472, 26613, 25471, 25997, 25710, 25367, 25020, 
    24562, 24021,
  24450, 24308, 25689, 25995, 26016, 25280, 24057, 23219, 22703, 22655, 
    22829, 23278, 24013, 25472, 26610, 25527, 25848, 25573, 25367, 25063, 
    24441, 24075,
  24593, 24460, 25798, 26022, 26001, 25305, 24019, 23213, 22727, 22624, 
    22900, 23319, 24047, 25376, 26194, 25571, 25804, 25479, 25325, 24957, 
    24492, 24115,
  24719, 24598, 25925, 26129, 26071, 25308, 24043, 23183, 22774, 22658, 
    22943, 23344, 24235, 25204, 26720, 25741, 26078, 25703, 25367, 24951, 
    24517, 24028,
  24792, 24696, 26016, 26181, 26097, 25316, 24019, 23178, 22735, 22583, 
    22926, 23347, 24264, 25430, 26420, 25875, 26078, 25732, 25353, 25020, 
    24479, 23987,
  24776, 24715, 25862, 26149, 26037, 25266, 24009, 23189, 22741, 22644, 
    22909, 23327, 24131, 25306, 26662, 25689, 26110, 25776, 25381, 24989, 
    24460, 24121,
  24641, 24617, 25837, 26041, 25997, 25246, 24005, 23162, 22735, 22652, 
    22900, 23296, 24220, 25418, 26572, 25591, 26159, 25782, 25374, 25032, 
    24485, 24055,
  24374, 24384, 25842, 26057, 26028, 25232, 23988, 23198, 22741, 22661, 
    22900, 23274, 24230, 25358, 26279, 25624, 26396, 26029, 25581, 25038, 
    24543, 24048,
  23976, 24019, 25781, 26087, 26014, 25204, 24026, 23234, 22718, 22658, 
    22906, 23350, 23936, 25283, 26384, 25521, 26601, 26245, 25719, 25169, 
    24555, 24068,
  23444, 23517, 25517, 25904, 25907, 25249, 24009, 23181, 22774, 22658, 
    22838, 23393, 24114, 25430, 26653, 25162, 26540, 26382, 25795, 25213, 
    24505, 24108,
  22748, 22831, 25154, 25681, 25865, 25243, 23971, 23172, 22759, 22656, 
    22886, 23307, 24116, 25390, 26388, 24908, 26490, 26462, 25871, 25294, 
    24632, 24162,
  21833, 21906, 24728, 25436, 25757, 25224, 23981, 23178, 22751, 22690, 
    22978, 23378, 24304, 25423, 26539, 24496, 26365, 26513, 25954, 25350, 
    24581, 24115,
  20696, 20760, 23957, 25051, 25610, 25112, 23954, 23213, 22739, 22616, 
    22906, 23299, 24371, 25337, 26231, 23900, 26310, 26628, 26051, 25518, 
    24760, 24196,
  19456, 19525, 23057, 24404, 25304, 25008, 23943, 23184, 22768, 22696, 
    22935, 23350, 24126, 25402, 26682, 22942, 25829, 26614, 26169, 25599, 
    24792, 24229,
  18343, 18421, 22244, 23947, 25115, 24972, 23905, 23140, 22757, 22736, 
    22949, 23373, 24161, 25281, 26444, 22051, 25300, 26635, 26203, 25660, 
    24798, 24129,
  17574, 17649, 21985, 23708, 25015, 24972, 23909, 23164, 22748, 22708, 
    22970, 23409, 24196, 25540, 26425, 21727, 25332, 26614, 26224, 25612, 
    24868, 24310,
  17246, 17302, 21960, 23727, 25001, 24893, 23902, 23158, 22751, 22725, 
    22893, 23338, 24068, 25384, 26826, 21713, 25163, 26563, 26321, 25749, 
    25047, 24304,
  17318, 17361, 22105, 23732, 24993, 24868, 23892, 23158, 22757, 22742, 
    22970, 23328, 24250, 25466, 26529, 21702, 25107, 26571, 26328, 25835, 
    25054, 24444,
  17692, 17741, 22120, 23724, 24984, 24914, 23864, 23173, 22757, 22760, 
    22890, 23439, 24320, 25533, 26379, 21735, 24964, 26585, 26349, 25892, 
    25111, 24424,
  18262, 18342, 22310, 23873, 24987, 24824, 23829, 23102, 22816, 22803, 
    22976, 23443, 24231, 25295, 26326, 21940, 24996, 26643, 26342, 25929, 
    25143, 24538,
  18923, 19037, 22790, 24142, 25073, 24860, 23805, 23097, 22822, 22723, 
    22876, 23389, 24044, 25179, 26663, 22400, 25133, 26607, 26384, 25917, 
    25207, 24418,
  19539, 19677, 23345, 24462, 25170, 24832, 23812, 23109, 22773, 22706, 
    22947, 23380, 24202, 25445, 26195, 23040, 25500, 26607, 26342, 25917, 
    25213, 24619,
  19959, 20120, 23705, 24696, 25257, 24830, 23802, 23100, 22790, 22781, 
    22936, 23415, 24111, 25247, 26612, 23513, 25687, 26499, 26342, 25849, 
    25277, 24592,
  20078, 20284, 23827, 24742, 25288, 24841, 23743, 23112, 22761, 22795, 
    22985, 23388, 24242, 25417, 26656, 23624, 25719, 26629, 26322, 25910, 
    25188, 24599,
  19894, 20159, 23672, 24710, 25251, 24805, 23750, 23106, 22802, 22778, 
    22991, 23466, 24353, 25664, 26876, 23417, 25532, 26629, 26404, 25918, 
    25259, 24707,
  19492, 19791, 23338, 24490, 25208, 24799, 23715, 23091, 22811, 22813, 
    22963, 23357, 24222, 25364, 26579, 23049, 25314, 26529, 26335, 25812, 
    25246, 24673,
  18992, 19268, 23034, 24301, 25074, 24760, 23715, 23110, 22808, 22839, 
    23029, 23614, 24336, 25569, 26438, 22612, 25202, 26529, 26343, 25843, 
    25252, 24740,
  18473, 18692, 22682, 24105, 25022, 24730, 23678, 23074, 22821, 22854, 
    22926, 23441, 24348, 25480, 26804, 22084, 24922, 26515, 26232, 25751, 
    25164, 24613,
  17955, 18137, 22426, 24019, 24983, 24705, 23671, 23092, 22789, 22811, 
    22992, 23526, 24383, 25544, 26610, 21811, 24960, 26443, 26192, 25745, 
    25100, 24600,
  17433, 17618, 22214, 23847, 24954, 24671, 23678, 23099, 22797, 22828, 
    23101, 23551, 24334, 25567, 26656, 21529, 24804, 26464, 26178, 25676, 
    25183, 24601,
  16923, 17120, 22039, 23799, 24897, 24576, 23592, 23043, 22806, 22854, 
    23047, 23468, 24396, 25432, 26641, 21361, 24774, 26450, 26116, 25676, 
    25139, 24594,
  16485, 16658, 21958, 23772, 24902, 24585, 23609, 23061, 22859, 22857, 
    23015, 23420, 24324, 25534, 26606, 21308, 24998, 26450, 26178, 25682, 
    25101, 24608,
  16198, 16318, 22077, 23888, 24948, 24568, 23602, 23064, 22857, 22843, 
    23033, 23597, 24359, 25700, 26460, 21355, 25023, 26428, 26206, 25739, 
    25158, 24688,
  16155, 16236, 22105, 23915, 24909, 24526, 23578, 22996, 22837, 22852, 
    23028, 23491, 24411, 25672, 26562, 21432, 25091, 26407, 26157, 25714, 
    25222, 24796,
  16472, 16557, 22296, 23982, 24957, 24526, 23578, 23023, 22869, 22861, 
    23127, 23474, 24456, 25719, 26695, 21529, 25198, 26429, 26144, 25739, 
    25197, 24682,
  17259, 17356, 22658, 24225, 25006, 24490, 23547, 23070, 22834, 22904, 
    23045, 23527, 24399, 25488, 26587, 21852, 25335, 26457, 26131, 25751, 
    25032, 24616,
  18503, 18563, 23355, 24524, 25052, 24479, 23478, 23000, 22814, 22888, 
    22960, 23543, 24432, 25691, 26466, 22565, 25565, 26435, 26089, 25622, 
    24969, 24348,
  19971, 19941, 24215, 24943, 25101, 24426, 23478, 22997, 22861, 22859, 
    23082, 23619, 24311, 25626, 26918, 23509, 25951, 26466, 26110, 25684, 
    25007, 24469,
  21290, 21181, 24749, 25231, 25158, 24415, 23423, 23000, 22794, 22808, 
    23068, 23660, 24405, 25766, 26860, 24159, 26150, 26415, 26104, 25653, 
    25065, 24583,
  22189, 22068, 24965, 25269, 25199, 24336, 23385, 22969, 22862, 22886, 
    23029, 23663, 24578, 25787, 26835, 24270, 25907, 26401, 26082, 25579, 
    24976, 24450,
  22685, 22609, 24808, 25245, 25096, 24292, 23368, 22945, 22847, 22886, 
    23035, 23615, 24696, 25954, 26810, 23915, 25901, 26279, 26007, 25567, 
    25027, 24524,
  23005, 22981, 24839, 25240, 25096, 24256, 23375, 22987, 22827, 22943, 
    23124, 23688, 24529, 25803, 27007, 23775, 25778, 26357, 26001, 25530, 
    24964, 24450,
  23329, 23322, 25285, 25493, 25145, 24264, 23341, 22975, 22862, 22964, 
    23141, 23615, 24689, 25759, 26848, 24562, 26381, 26401, 26035, 25537, 
    25009, 24638,
  23616, 23598, 25812, 25706, 25211, 24189, 23303, 22940, 22851, 22898, 
    23190, 23593, 24650, 25897, 26829, 25488, 26835, 26445, 25988, 25537, 
    24996, 24458,
  23691, 23677, 25903, 25760, 25176, 24184, 23234, 22908, 22854, 22893, 
    23215, 23684, 24577, 25926, 26726, 25666, 26704, 26323, 25981, 25500, 
    24946, 24365,
  23439, 23457, 25660, 25644, 25062, 24100, 23238, 22920, 22851, 22916, 
    23125, 23700, 24761, 25890, 27204, 25454, 26568, 26309, 25947, 25500, 
    24806, 24258,
  22881, 22892, 25366, 25453, 24991, 24049, 23210, 22914, 22863, 22985, 
    23301, 23783, 24703, 26109, 26846, 24773, 26413, 26244, 25871, 25432, 
    24845, 24232,
  22140, 22028, 25027, 25295, 24894, 23988, 23158, 22879, 22858, 22939, 
    23205, 23807, 24723, 26057, 27384, 23538, 26176, 26251, 25837, 25370, 
    24889, 24339,
  21469, 21163, 24961, 25230, 24845, 23913, 23110, 22909, 22864, 23022, 
    23142, 23880, 24841, 26391, 27040, 23130, 26132, 26100, 25734, 25265, 
    24725, 24192,
  21193, 20789, 25174, 25300, 24762, 23837, 23078, 22892, 22864, 23043, 
    23276, 23784, 24918, 25941, 26596, 23459, 26109, 26035, 25569, 25147, 
    24483, 24032,
  28593, 28516, 27844, 27118, 25760, 24108, 22722, 22183, 22085, 22499, 
    23039, 23629, 24590, 25875, 26601, 28588, 28907, 27966, 27374, 26562, 
    25407, 24408,
  28573, 28511, 27913, 27201, 25914, 24245, 22798, 22201, 22099, 22504, 
    22885, 23621, 24550, 25854, 26734, 28582, 28801, 27865, 27250, 26431, 
    25368, 24362,
  28527, 28497, 27844, 27215, 25945, 24352, 22860, 22233, 22151, 22573, 
    22881, 23633, 24530, 25891, 26887, 28532, 28676, 27706, 27104, 26382, 
    25279, 24228,
  28470, 28476, 27810, 27298, 26066, 24452, 22929, 22324, 22116, 22478, 
    22913, 23534, 24549, 25621, 26671, 28541, 28589, 27612, 26954, 26107, 
    25113, 24054,
  28404, 28436, 27913, 27204, 26148, 24522, 23009, 22356, 22154, 22515, 
    22915, 23493, 24495, 25729, 26526, 28518, 28501, 27532, 26829, 26015, 
    24897, 23973,
  28318, 28360, 27829, 27263, 26197, 24631, 23054, 22394, 22200, 22483, 
    22818, 23541, 24520, 25523, 26920, 28443, 28409, 27482, 26788, 25951, 
    24884, 24020,
  28199, 28231, 27801, 27231, 26217, 24692, 23137, 22435, 22165, 22457, 
    22849, 23523, 24554, 25784, 26601, 28367, 28341, 27179, 26553, 25766, 
    24827, 23979,
  28034, 28047, 27750, 27268, 26254, 24762, 23216, 22488, 22191, 22485, 
    22803, 23480, 24278, 25700, 26816, 28219, 28041, 26804, 26084, 25374, 
    24490, 23912,
  27831, 27828, 27563, 27157, 26201, 24762, 23241, 22491, 22246, 22516, 
    22920, 23444, 24410, 25595, 26734, 28082, 27804, 26609, 25925, 25275, 
    24508, 23905,
  27627, 27613, 27387, 27039, 26179, 24852, 23341, 22564, 22245, 22482, 
    22840, 23454, 24457, 25490, 26615, 27700, 27469, 26292, 25712, 25188, 
    24521, 24025,
  27471, 27444, 27116, 26835, 26104, 24871, 23327, 22584, 22269, 22464, 
    22930, 23542, 24531, 25452, 26959, 27160, 26741, 26003, 25587, 25144, 
    24514, 24038,
  27399, 27347, 26896, 26668, 26010, 24871, 23375, 22601, 22280, 22470, 
    22867, 23474, 24292, 25557, 26663, 26700, 25676, 25577, 25401, 24988, 
    24393, 23817,
  27419, 27332, 26923, 26681, 26028, 24916, 23465, 22622, 22318, 22438, 
    22902, 23400, 24471, 25464, 26513, 26539, 24986, 25159, 25084, 24882, 
    24304, 23864,
  27493, 27381, 26997, 26778, 26122, 24870, 23496, 22672, 22359, 22520, 
    22870, 23440, 24409, 25618, 26726, 26701, 25123, 25202, 25118, 24938, 
    24361, 23917,
  27553, 27442, 27132, 26829, 26196, 24960, 23496, 22698, 22311, 22560, 
    22867, 23410, 24337, 25436, 26554, 26843, 25888, 25519, 25331, 24938, 
    24341, 23970,
  27538, 27445, 27101, 26875, 26247, 25007, 23603, 22736, 22329, 22443, 
    22852, 23397, 24327, 25303, 26687, 26904, 25763, 25447, 25324, 24913, 
    24360, 23829,
  27445, 27360, 27189, 26882, 26284, 25052, 23610, 22792, 22361, 22517, 
    22889, 23419, 24300, 25526, 26498, 26953, 25800, 25476, 25227, 24900, 
    24226, 23809,
  27313, 27222, 27047, 26885, 26273, 25077, 23669, 22780, 22404, 22488, 
    22835, 23436, 24280, 25291, 26415, 27145, 26578, 25850, 25427, 24980, 
    24359, 23701,
  27198, 27103, 26948, 26776, 26284, 25147, 23690, 22818, 22416, 22537, 
    22868, 23510, 24280, 25622, 26493, 27165, 26995, 26175, 25647, 25049, 
    24339, 23855,
  27135, 27048, 26892, 26818, 26275, 25166, 23738, 22873, 22465, 22464, 
    22808, 23452, 24300, 25516, 26321, 27185, 27175, 26290, 25716, 25054, 
    24320, 23754,
  27117, 27051, 27037, 26867, 26316, 25183, 23738, 22894, 22474, 22542, 
    22876, 23332, 24295, 25390, 26535, 27321, 26970, 26160, 25606, 24961, 
    24288, 23754,
  27113, 27079, 27201, 26957, 26289, 25147, 23779, 22941, 22464, 22518, 
    22811, 23461, 24252, 25320, 26720, 27413, 26839, 26066, 25585, 24960, 
    24383, 23687,
  27111, 27107, 27196, 26917, 26347, 25230, 23804, 22982, 22476, 22515, 
    22862, 23380, 24213, 25279, 26676, 27432, 26764, 26079, 25591, 24972, 
    24345, 23706,
  27140, 27127, 27123, 26920, 26347, 25239, 23838, 22976, 22485, 22544, 
    22867, 23400, 24207, 25437, 26426, 27434, 26726, 26044, 25619, 25097, 
    24408, 23740,
  27223, 27156, 27176, 26982, 26375, 25275, 23855, 22987, 22522, 22523, 
    22913, 23364, 24247, 25411, 26679, 27531, 26901, 26123, 25722, 25183, 
    24459, 23820,
  27333, 27218, 27341, 27071, 26447, 25286, 23900, 23019, 22552, 22538, 
    22858, 23422, 24249, 25406, 26339, 27612, 27169, 26360, 25819, 25258, 
    24510, 23986,
  27412, 27311, 27260, 27051, 26407, 25339, 23896, 23010, 22572, 22537, 
    22775, 23356, 24244, 25169, 26504, 27509, 27206, 26354, 25929, 25277, 
    24484, 23866,
  27423, 27391, 27226, 26925, 26378, 25297, 23900, 23001, 22545, 22531, 
    22830, 23455, 24239, 25434, 26543, 27392, 27013, 26303, 25832, 25270, 
    24579, 23999,
  27371, 27395, 27117, 26919, 26315, 25286, 23910, 23066, 22577, 22511, 
    22835, 23371, 24270, 25346, 26194, 27307, 26913, 26245, 25797, 25276, 
    24521, 23972,
  27255, 27292, 27092, 26925, 26282, 25314, 23927, 23066, 22545, 22551, 
    22866, 23409, 24086, 25299, 26414, 27254, 26820, 26216, 25742, 25195, 
    24464, 23992,
  27055, 27079, 27059, 26832, 26289, 25224, 23962, 23057, 22554, 22562, 
    22843, 23282, 24122, 25368, 26443, 27228, 26720, 26216, 25790, 25288, 
    24610, 23851,
  26745, 26761, 27009, 26782, 26266, 25313, 23934, 23066, 22618, 22539, 
    22892, 23357, 24248, 25387, 26297, 27182, 26826, 26223, 25741, 25220, 
    24463, 23958,
  26330, 26343, 26838, 26707, 26220, 25249, 23923, 23071, 22609, 22530, 
    22880, 23330, 24203, 25312, 26104, 27142, 26795, 26135, 25728, 25288, 
    24546, 23965,
  25857, 25861, 26643, 26566, 26179, 25280, 23975, 23095, 22556, 22530, 
    22888, 23360, 24322, 25445, 26416, 27010, 26539, 26129, 25769, 25350, 
    24654, 24038,
  25395, 25401, 26470, 26467, 26131, 25229, 23930, 23121, 22588, 22564, 
    22905, 23314, 24287, 25338, 26079, 26871, 26545, 26013, 25657, 25312, 
    24629, 24065,
  25016, 25055, 26307, 26389, 26045, 25201, 23982, 23095, 22612, 22622, 
    22871, 23266, 24247, 25219, 26329, 26765, 26432, 25956, 25589, 25132, 
    24609, 24005,
  24787, 24867, 26135, 26254, 26016, 25237, 23968, 23121, 22661, 22509, 
    22794, 23283, 24161, 25312, 26525, 26626, 26332, 25904, 25562, 25150, 
    24571, 23984,
  24747, 24814, 26059, 26235, 25994, 25218, 23996, 23136, 22635, 22636, 
    22928, 23331, 24161, 25331, 26310, 26476, 26271, 25775, 25499, 25156, 
    24565, 24104,
  24854, 24840, 26153, 26249, 26025, 25265, 23989, 23171, 22679, 22621, 
    22867, 23326, 24099, 25382, 26365, 26250, 26121, 25760, 25492, 25132, 
    24558, 24024,
  24983, 24875, 26160, 26229, 26057, 25263, 24010, 23159, 22660, 22569, 
    22873, 23288, 24087, 25368, 26840, 26135, 25853, 25753, 25485, 25225, 
    24679, 24084,
  25004, 24848, 26064, 26275, 26071, 25218, 24006, 23189, 22707, 22615, 
    22796, 23361, 24163, 25200, 26201, 26239, 26151, 25818, 25499, 25125, 
    24551, 23997,
  24874, 24715, 25942, 26176, 26037, 25310, 24041, 23159, 22678, 22601, 
    22873, 23278, 24123, 25216, 26748, 26110, 26532, 25954, 25513, 25144, 
    24513, 24077,
  24654, 24503, 25798, 26063, 26034, 25296, 24034, 23230, 22757, 22578, 
    22856, 23313, 24207, 25179, 26263, 25904, 26626, 25984, 25506, 25144, 
    24526, 23944,
  24453, 24307, 25813, 26084, 25996, 25290, 23999, 23171, 22704, 22652, 
    22987, 23343, 24047, 25160, 26560, 25885, 26619, 25991, 25513, 25031, 
    24474, 23950,
  24351, 24211, 25773, 26062, 25988, 25257, 23985, 23144, 22748, 22592, 
    22807, 23313, 24089, 25261, 26178, 25771, 26563, 25984, 25568, 25019, 
    24526, 23983,
  24358, 24224, 25653, 25954, 25999, 25226, 24023, 23165, 22730, 22644, 
    22801, 23333, 24387, 25160, 26504, 25504, 26451, 26004, 25623, 25119, 
    24551, 24050,
  24431, 24302, 25585, 25954, 25956, 25254, 24003, 23165, 22733, 22618, 
    22910, 23321, 24237, 25268, 26651, 25396, 26270, 25932, 25506, 25087, 
    24462, 23903,
  24523, 24398, 25726, 25976, 26019, 25310, 24003, 23236, 22777, 22658, 
    22787, 23346, 24077, 25361, 26420, 25451, 26051, 25781, 25416, 25057, 
    24519, 24017,
  24612, 24500, 25793, 26014, 25988, 25248, 24020, 23182, 22748, 22621, 
    22836, 23316, 24128, 25407, 26029, 25518, 25785, 25485, 25278, 24888, 
    24373, 23930,
  24693, 24604, 25945, 26165, 26082, 25271, 23995, 23191, 22751, 22658, 
    22779, 23336, 24146, 25249, 26445, 25704, 25710, 25312, 25091, 24777, 
    24411, 23943,
  24754, 24695, 26018, 26203, 26068, 25274, 23975, 23183, 22739, 22666, 
    22881, 23369, 24190, 25358, 26357, 25851, 26345, 25796, 25374, 24938, 
    24544, 23896,
  24768, 24739, 26095, 26207, 26101, 25301, 23992, 23188, 22745, 22649, 
    22899, 23397, 24079, 25249, 26316, 25876, 26464, 25825, 25443, 24982, 
    24455, 23943,
  24701, 24694, 25982, 26159, 26056, 25262, 24023, 23206, 22748, 22669, 
    22839, 23267, 24170, 25137, 26579, 25782, 26451, 25984, 25519, 24969, 
    24443, 23944,
  24524, 24537, 25907, 26157, 26062, 25220, 24006, 23221, 22775, 22647, 
    22930, 23336, 24168, 25268, 26549, 25760, 26588, 26085, 25651, 25088, 
    24500, 24010,
  24216, 24258, 25788, 26098, 26037, 25240, 24023, 23206, 22757, 22701, 
    22845, 23359, 24222, 25342, 26504, 25671, 26682, 26222, 25713, 25162, 
    24545, 24037,
  23745, 23826, 25562, 25966, 25968, 25223, 24020, 23218, 22719, 22687, 
    22850, 23293, 24183, 25333, 26348, 25375, 26676, 26403, 25857, 25299, 
    24557, 24057,
  23051, 23158, 25410, 25831, 25891, 25204, 23971, 23195, 22784, 22613, 
    22947, 23309, 24242, 25401, 26353, 25108, 26620, 26562, 25926, 25411, 
    24647, 24131,
  22056, 22175, 24926, 25511, 25770, 25167, 23982, 23177, 22775, 22699, 
    22913, 23369, 24099, 25389, 26479, 24648, 26532, 26670, 26072, 25380, 
    24724, 24051,
  20749, 20887, 23812, 24862, 25504, 25072, 23975, 23183, 22766, 22664, 
    22911, 23372, 24210, 25338, 26646, 23465, 25878, 26641, 26251, 25604, 
    24895, 24185,
  19270, 19446, 22499, 24027, 25158, 24971, 23916, 23201, 22781, 22748, 
    22933, 23410, 24047, 25233, 26644, 21955, 25194, 26591, 26238, 25648, 
    24806, 24272,
  17895, 18109, 21855, 23648, 24995, 24962, 23926, 23166, 22807, 22730, 
    22971, 23362, 24319, 25235, 26494, 21279, 25119, 26569, 26224, 25648, 
    24889, 24111,
  16913, 17135, 21949, 23691, 24995, 24921, 23906, 23136, 22831, 22682, 
    22919, 23441, 24193, 25443, 26814, 21582, 25412, 26576, 26287, 25673, 
    24941, 24326,
  16484, 16684, 22094, 23702, 24966, 24918, 23902, 23184, 22790, 22785, 
    22874, 23398, 24344, 25401, 26789, 21788, 25430, 26554, 26287, 25723, 
    24953, 24433,
  16604, 16770, 22038, 23715, 24981, 24907, 23868, 23204, 22802, 22791, 
    22925, 23411, 24152, 25573, 26646, 21709, 25219, 26606, 26404, 25829, 
    24966, 24399,
  17148, 17290, 22054, 23724, 24978, 24857, 23843, 23178, 22776, 22763, 
    23034, 23416, 24374, 25264, 26654, 21611, 24957, 26541, 26307, 25879, 
    25056, 24333,
  17947, 18076, 22343, 23950, 25012, 24826, 23837, 23134, 22759, 22777, 
    22954, 23376, 24150, 25529, 26646, 21878, 25007, 26570, 26391, 25817, 
    25094, 24427,
  18822, 18946, 22923, 24230, 25119, 24893, 23827, 23116, 22802, 22821, 
    23060, 23434, 24307, 25467, 26598, 22496, 25281, 26520, 26342, 25848, 
    25081, 24440,
  19601, 19731, 23519, 24561, 25213, 24834, 23830, 23190, 22826, 22778, 
    22966, 23404, 24275, 25383, 26613, 23128, 25593, 26628, 26343, 25885, 
    25075, 24427,
  20147, 20306, 23813, 24758, 25268, 24851, 23785, 23123, 22765, 22795, 
    22946, 23488, 24194, 25506, 26868, 23548, 25660, 26570, 26412, 25892, 
    25197, 24428,
  20392, 20609, 23773, 24747, 25310, 24815, 23796, 23096, 22800, 22801, 
    23001, 23414, 24375, 25523, 26501, 23545, 25643, 26614, 26350, 25898, 
    25177, 24642,
  20346, 20635, 23611, 24710, 25208, 24796, 23754, 23090, 22830, 22830, 
    23004, 23470, 24330, 25592, 26604, 23341, 25469, 26570, 26343, 25849, 
    25241, 24541,
  20079, 20413, 23449, 24583, 25222, 24756, 23727, 23097, 22789, 22836, 
    23024, 23503, 24392, 25542, 26760, 23051, 25264, 26556, 26301, 25762, 
    25159, 24562,
  19675, 19997, 23350, 24478, 25153, 24774, 23744, 23091, 22809, 22759, 
    23084, 23451, 24311, 25756, 26717, 22906, 25288, 26506, 26274, 25737, 
    25184, 24589,
  19195, 19464, 23165, 24347, 25119, 24734, 23724, 23088, 22865, 22865, 
    23044, 23456, 24254, 25574, 26529, 22596, 25226, 26463, 26212, 25694, 
    25038, 24602,
  18655, 18883, 22889, 24307, 25099, 24704, 23685, 23085, 22822, 22820, 
    23064, 23420, 24467, 25465, 26487, 22337, 25127, 26419, 26129, 25706, 
    25007, 24556,
  18054, 18276, 22725, 24154, 25022, 24656, 23651, 23068, 22822, 22928, 
    23048, 23489, 24390, 25817, 26645, 22052, 25108, 26434, 26137, 25620, 
    25102, 24489,
  17416, 17641, 22408, 24019, 24931, 24634, 23651, 23107, 22831, 22863, 
    23082, 23484, 24341, 25593, 27098, 21731, 24953, 26348, 26060, 25545, 
    24982, 24523,
  16815, 17014, 22206, 23922, 24899, 24595, 23606, 23030, 22849, 22869, 
    23148, 23553, 24366, 25665, 26732, 21497, 24935, 26449, 26129, 25695, 
    25052, 24470,
  16366, 16515, 22133, 23844, 24954, 24553, 23578, 23122, 22858, 22886, 
    23068, 23462, 24465, 25678, 26762, 21393, 25003, 26413, 26185, 25751, 
    25110, 24711,
  16216, 16329, 22219, 23942, 24929, 24592, 23589, 23081, 22899, 22887, 
    23145, 23587, 24470, 25510, 26929, 21456, 25122, 26500, 26151, 25776, 
    25142, 24597,
  16523, 16636, 22374, 24025, 24989, 24542, 23572, 23084, 22873, 22967, 
    23112, 23579, 24335, 25720, 26825, 21665, 25215, 26457, 26172, 25838, 
    25206, 24651,
  17390, 17506, 22774, 24243, 24992, 24506, 23531, 23026, 22870, 22910, 
    23001, 23592, 24574, 25825, 27176, 22068, 25464, 26399, 26069, 25651, 
    24977, 24484,
  18748, 18823, 23484, 24553, 25078, 24469, 23489, 23043, 22838, 22936, 
    23030, 23574, 24454, 25687, 27092, 22854, 25838, 26370, 26000, 25547, 
    24933, 24331,
  20298, 20293, 24308, 24997, 25155, 24447, 23496, 23032, 22871, 22954, 
    23084, 23666, 24513, 25536, 26851, 23804, 26079, 26378, 26021, 25566, 
    24952, 24371,
  21631, 21561, 24860, 25247, 25207, 24445, 23479, 22985, 22827, 22868, 
    23207, 23542, 24535, 26069, 27038, 24356, 26137, 26371, 26021, 25560, 
    25054, 24485,
  22480, 22402, 25000, 25328, 25204, 24353, 23455, 23000, 22851, 22960, 
    23127, 23649, 24447, 25790, 26626, 24373, 26044, 26335, 25939, 25504, 
    24991, 24392,
  22882, 22841, 24944, 25258, 25181, 24322, 23403, 22997, 22860, 22977, 
    23136, 23589, 24561, 25795, 26810, 24096, 26044, 26220, 25856, 25467, 
    24851, 24359,
  23094, 23087, 24937, 25296, 25150, 24305, 23393, 22968, 22901, 22940, 
    23173, 23677, 24630, 25842, 26925, 23970, 25926, 26204, 25794, 25362, 
    24794, 24239,
  23328, 23321, 25277, 25503, 25204, 24294, 23331, 22968, 22863, 22926, 
    23168, 23705, 24689, 25929, 26821, 24625, 26274, 26213, 25870, 25374, 
    24763, 24326,
  23579, 23557, 25740, 25735, 25230, 24239, 23307, 22978, 22905, 22938, 
    23211, 23782, 24643, 25793, 27157, 25549, 26729, 26307, 25829, 25418, 
    24782, 24367,
  23698, 23688, 25869, 25762, 25147, 24155, 23283, 22998, 22858, 22976, 
    23200, 23739, 24700, 26144, 26854, 25735, 26704, 26250, 25801, 25369, 
    24783, 24253,
  23562, 23596, 25682, 25606, 25073, 24113, 23231, 22963, 22899, 22979, 
    23240, 23769, 24786, 26124, 27206, 25339, 26443, 26235, 25837, 25369, 
    24770, 24160,
  23137, 23175, 25376, 25413, 25008, 24049, 23210, 22928, 22882, 23034, 
    23189, 23777, 24818, 25828, 26959, 24744, 26368, 26257, 25844, 25381, 
    24783, 24288,
  22490, 22418, 25067, 25273, 24888, 24007, 23158, 22946, 22900, 22985, 
    23198, 23929, 24764, 26212, 27192, 23682, 26219, 26228, 25837, 25407, 
    24796, 24308,
  21855, 21603, 25006, 25248, 24831, 23873, 23110, 22937, 22903, 22971, 
    23269, 23874, 24720, 26115, 27001, 23375, 26231, 26091, 25769, 25333, 
    24720, 24188,
  21584, 21242, 25192, 25268, 24762, 23806, 23093, 22946, 22871, 23020, 
    23204, 23829, 24752, 26084, 27232, 23628, 26182, 25912, 25534, 25091, 
    24397, 23961 ;
}
