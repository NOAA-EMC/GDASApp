netcdf rads_adt_3a_2021182 {
dimensions:
	time = UNLIMITED ; // (11 currently)
variables:
	int adt_egm2008(time) ;
		adt_egm2008:_FillValue = 2147483647 ;
		adt_egm2008:long_name = "absolute dynamic topography (EGM2008)" ;
		adt_egm2008:standard_name = "absolute_dynamic_topography_egm2008" ;
		adt_egm2008:units = "m" ;
		adt_egm2008:scale_factor = 0.0001 ;
		adt_egm2008:coordinates = "lon lat" ;
	int adt_xgm2016(time) ;
		adt_xgm2016:_FillValue = 2147483647 ;
		adt_xgm2016:long_name = "absolute dynamic topography (XGM2016)" ;
		adt_xgm2016:standard_name = "absolute_dynamic_topography_xgm2016" ;
		adt_xgm2016:units = "m" ;
		adt_xgm2016:scale_factor = 0.0001 ;
		adt_xgm2016:coordinates = "lon lat" ;
	int cycle(time) ;
		cycle:_FillValue = 2147483647 ;
		cycle:long_name = "cycle number" ;
		cycle:field = 9905s ;
	int lat(time) ;
		lat:_FillValue = 2147483647 ;
		lat:long_name = "latitude" ;
		lat:standard_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:scale_factor = 1.e-06 ;
		lat:field = 201s ;
		lat:comment = "Positive latitude is North latitude, negative latitude is South latitude" ;
	int lon(time) ;
		lon:_FillValue = 2147483647 ;
		lon:long_name = "longitude" ;
		lon:standard_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:scale_factor = 1.e-06 ;
		lon:field = 301s ;
		lon:comment = "East longitude relative to Greenwich meridian" ;
	int pass(time) ;
		pass:_FillValue = 2147483647 ;
		pass:long_name = "pass number" ;
		pass:field = 9906s ;
	short sla(time) ;
		sla:_FillValue = 32767s ;
		sla:long_name = "sea level anomaly" ;
		sla:standard_name = "sea_surface_height_above_sea_level" ;
		sla:units = "m" ;
		sla:quality_flag = "swh sig0 range_rms range_numval flags swh_rms sig0_rms" ;
		sla:scale_factor = 0.0001 ;
		sla:coordinates = "lon lat" ;
		sla:field = 0s ;
		sla:comment = "Sea level determined from satellite altitude - range - all altimetric corrections" ;
	double time_dtg(time) ;
		time_dtg:long_name = "time_dtg" ;
		time_dtg:standard_name = "time_dtg" ;
		time_dtg:units = "yyyymmddhhmmss" ;
		time_dtg:coordinates = "lon lat" ;
		time_dtg:comment = "UTC time formatted as yyyymmddhhmmss" ;
	double time_mjd(time) ;
		time_mjd:long_name = "Modified Julian Days" ;
		time_mjd:standard_name = "time" ;
		time_mjd:units = "days since 1858-11-17 00:00:00 UTC" ;
		time_mjd:field = 105s ;
		time_mjd:comment = "UTC time of measurement expressed in Modified Julian Days" ;

// global attributes:
		:Conventions = "CF-1.7" ;
		:title = "RADS 4 pass file" ;
		:institution = "EUMETSAT / NOAA / TU Delft" ;
		:source = "radar altimeter" ;
		:references = "RADS Data Manual, Version 4.2 or later" ;
		:featureType = "trajectory" ;
		:ellipsoid = "TOPEX" ;
		:ellipsoid_axis = 6378136.3 ;
		:ellipsoid_flattening = 0.00335281317789691 ;
		:filename = "rads_adt_3a_2021182.nc" ;
		:mission_name = "SNTNL-3A" ;
		:mission_phase = "a" ;
		:log01 = "2021-07-02 | /Users/rads/bin/rads2nc --ymd=20210701000000,20210702000000 -C1,1000 -S3a -Vsla,adt_egm2008,adt_xgm2016,time_mjd,time_dtg,lon,lat,cycle,pass -X/Users/rads/cron/xgm2016 -X/Users/rads/cron/adt -X/Users/rads/cron/time_dtg -o/Users/rads/adt/2021/182/rads_adt_3a_2021182.nc: RAW data from" ;
		:history = "Mon Sep 25 17:01:31 2023: ncks -d time,0,10 rads_adt_3a_2021182.nc rads_adt_3a_2021182.ncn\n",
			"2021-07-02 21:11:15 : /Users/rads/bin/rads2nc --ymd=20210701000000,20210702000000 -C1,1000 -S3a -Vsla,adt_egm2008,adt_xgm2016,time_mjd,time_dtg,lon,lat,cycle,pass -X/Users/rads/cron/xgm2016 -X/Users/rads/cron/adt -X/Users/rads/cron/time_dtg -o/Users/rads/adt/2021/182/rads_adt_3a_2021182.nc" ;
		:NCO = "netCDF Operators version 5.0.6 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco)" ;
data:

 adt_egm2008 = -4374, -3849, -3832, -3530, -3149, -2888, -2611, -2423, -2116, 
    -2011, -2170 ;

 adt_xgm2016 = -4617, -4012, -3779, -3212, -2781, -2466, -2048, -2067, -1971, 
    -2110, -2327 ;

 cycle = 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73 ;

 lat = 48396720, 48454663, 48512601, 48570535, 48628465, 48686391, 48744313, 
    48802230, 48860143, 48918052, 48975957 ;

 lon = -39706628, -39730940, -39755297, -39779700, -39804149, -39828645, 
    -39853187, -39877776, -39902412, -39927095, -39951826 ;

 pass = 545, 545, 545, 545, 545, 545, 545, 545, 545, 545, 545 ;

 sla = -3955, -3487, -3628, -3103, -2815, -2565, -2353, -2275, -1983, -1491, 
    -1688 ;

 time_dtg = 20210701000001, 20210701000002, 20210701000003, 20210701000004, 
    20210701000005, 20210701000006, 20210701000007, 20210701000008, 
    20210701000009, 20210701000010, 20210701000011 ;

 time_mjd = 59396.0000115741, 59396.0000231481, 59396.0000347222, 
    59396.0000462963, 59396.0000578704, 59396.0000694444, 59396.0000810185, 
    59396.0000925926, 59396.0001041667, 59396.0001157407, 59396.0001273148 ;
}
