netcdf sss_smos_1 {
dimensions:
	n_grid_points = 50 ;
variables:
	float A_card(n_grid_points) ;
		A_card:_FillValue = -999.f ;
	ubyte Coast_distance(n_grid_points) ;
		Coast_distance:_FillValue = 0UB ;
		Coast_distance:scale_factor = 20. ;
		Coast_distance:scale_offset = 0. ;
		string Coast_distance:_Unsigned = "true" ;
	uint Control_Flags_Acard(n_grid_points) ;
		Control_Flags_Acard:_FillValue = 0U ;
		Control_Flags_Acard:flag_masks = 2s, 4s, 8s, 16s, 32s, 64s, 128s, 256s, 512s, 1024s, 2048s, 4096s, 8192s, 16384s, -32768s, 0s, 0s, 0s, 0s, 0s, 0s, 0s, 0s, 0s, 0s, 0s, 0s, 0s, 0s ;
		Control_Flags_Acard:flag_values = 2s, 4s, 8s, 16s, 32s, 64s, 128s, 256s, 512s, 1024s, 2048s, 4096s, 8192s, 16384s, -32768s, 0s, 0s, 0s, 0s, 0s, 0s, 0s, 0s, 0s, 0s, 0s, 0s, 0s, 0s ;
		string Control_Flags_Acard:flag_meanings = "FG_CTRL_RANGE FG_CTRL_SIGMA FG_CTRL_CHI2 FG_CTRL_CHI2_P FG_CTRL_CONTAMINATED FG_CTRL_SUNGLINT FG_CTRL_MOONGLINT FG_CTRL_GAL_NOISE FG_CTRL_MIXED_SCENE FG_CTRL_REACH_MAXITER FG_CTRL_NUM_MEAS_MIN FG_CTRL_NUM_MEAS_LOW FG_CTRL_MANY_OUTLIERS FG_CTRL_MARQ FG_CTRL_ROUGHNESS FG_CTRL_FOAM FG_CTRL_ECMWF FG_CTRL_VALID FG_CTRL_NO_SURFACE FG_CTRL_RANGE_ACARD FG_CTRL_SIGMA_ACARD FG_CTRL_USED_FARATEC FG_CTRL_POOR_GEOPHYS FG_CTRL_POOR_RETRIEVAL FG_CTRL_SUSPECT_RFI FG_CTRL_RFI_PRONE_X FG_CTRL_RFI_PRONE_Y FG_CTRL_ADJUSTED_RA FG_CTRL_RETRIEV_FAIL" ;
		string Control_Flags_Acard:_Unsigned = "true" ;
	uint Control_Flags_anom(n_grid_points) ;
		Control_Flags_anom:_FillValue = 0U ;
		Control_Flags_anom:flag_masks = 2s, 4s, 8s, 16s, 32s, 64s, 128s, 256s, 512s, 1024s, 2048s, 4096s, 8192s, 16384s, -32768s, 0s, 0s, 0s, 0s, 0s, 0s, 0s, 0s, 0s, 0s, 0s, 0s, 0s, 0s ;
		Control_Flags_anom:flag_values = 2s, 4s, 8s, 16s, 32s, 64s, 128s, 256s, 512s, 1024s, 2048s, 4096s, 8192s, 16384s, -32768s, 0s, 0s, 0s, 0s, 0s, 0s, 0s, 0s, 0s, 0s, 0s, 0s, 0s, 0s ;
		string Control_Flags_anom:flag_meanings = "FG_CTRL_RANGE FG_CTRL_SIGMA FG_CTRL_CHI2 FG_CTRL_CHI2_P FG_CTRL_CONTAMINATED FG_CTRL_SUNGLINT FG_CTRL_MOONGLINT FG_CTRL_GAL_NOISE FG_CTRL_MIXED_SCENE FG_CTRL_REACH_MAXITER FG_CTRL_NUM_MEAS_MIN FG_CTRL_NUM_MEAS_LOW FG_CTRL_MANY_OUTLIERS FG_CTRL_MARQ FG_CTRL_ROUGHNESS FG_CTRL_FOAM FG_CTRL_ECMWF FG_CTRL_VALID FG_CTRL_NO_SURFACE FG_CTRL_RANGE_ACARD FG_CTRL_SIGMA_ACARD FG_CTRL_USED_FARATEC FG_CTRL_POOR_GEOPHYS FG_CTRL_POOR_RETRIEVAL FG_CTRL_SUSPECT_RFI FG_CTRL_RFI_PRONE_X FG_CTRL_RFI_PRONE_Y FG_CTRL_ADJUSTED_RA FG_CTRL_RETRIEV_FAIL" ;
		string Control_Flags_anom:_Unsigned = "true" ;
	uint Control_Flags_corr(n_grid_points) ;
		Control_Flags_corr:_FillValue = 0U ;
		Control_Flags_corr:flag_masks = 2s, 4s, 8s, 16s, 32s, 64s, 128s, 256s, 512s, 1024s, 2048s, 4096s, 8192s, 16384s, -32768s, 0s, 0s, 0s, 0s, 0s, 0s, 0s, 0s, 0s, 0s, 0s, 0s, 0s, 0s ;
		Control_Flags_corr:flag_values = 2s, 4s, 8s, 16s, 32s, 64s, 128s, 256s, 512s, 1024s, 2048s, 4096s, 8192s, 16384s, -32768s, 0s, 0s, 0s, 0s, 0s, 0s, 0s, 0s, 0s, 0s, 0s, 0s, 0s, 0s ;
		string Control_Flags_corr:flag_meanings = "FG_CTRL_RANGE FG_CTRL_SIGMA FG_CTRL_CHI2 FG_CTRL_CHI2_P FG_CTRL_CONTAMINATED FG_CTRL_SUNGLINT FG_CTRL_MOONGLINT FG_CTRL_GAL_NOISE FG_CTRL_MIXED_SCENE FG_CTRL_REACH_MAXITER FG_CTRL_NUM_MEAS_MIN FG_CTRL_NUM_MEAS_LOW FG_CTRL_MANY_OUTLIERS FG_CTRL_MARQ FG_CTRL_ROUGHNESS FG_CTRL_FOAM FG_CTRL_ECMWF FG_CTRL_VALID FG_CTRL_NO_SURFACE FG_CTRL_RANGE_ACARD FG_CTRL_SIGMA_ACARD FG_CTRL_USED_FARATEC FG_CTRL_POOR_GEOPHYS FG_CTRL_POOR_RETRIEVAL FG_CTRL_SUSPECT_RFI FG_CTRL_RFI_PRONE_X FG_CTRL_RFI_PRONE_Y FG_CTRL_ADJUSTED_RA FG_CTRL_RETRIEV_FAIL" ;
		string Control_Flags_corr:_Unsigned = "true" ;
	uint Control_Flags_uncorr(n_grid_points) ;
		Control_Flags_uncorr:_FillValue = 0U ;
		Control_Flags_uncorr:flag_masks = 2s, 4s, 8s, 16s, 32s, 64s, 128s, 256s, 512s, 1024s, 2048s, 4096s, 8192s, 16384s, -32768s, 0s, 0s, 0s, 0s, 0s, 0s, 0s, 0s, 0s, 0s, 0s, 0s, 0s, 0s ;
		Control_Flags_uncorr:flag_values = 2s, 4s, 8s, 16s, 32s, 64s, 128s, 256s, 512s, 1024s, 2048s, 4096s, 8192s, 16384s, -32768s, 0s, 0s, 0s, 0s, 0s, 0s, 0s, 0s, 0s, 0s, 0s, 0s, 0s, 0s ;
		string Control_Flags_uncorr:flag_meanings = "FG_CTRL_RANGE FG_CTRL_SIGMA FG_CTRL_CHI2 FG_CTRL_CHI2_P FG_CTRL_CONTAMINATED FG_CTRL_SUNGLINT FG_CTRL_MOONGLINT FG_CTRL_GAL_NOISE FG_CTRL_MIXED_SCENE FG_CTRL_REACH_MAXITER FG_CTRL_NUM_MEAS_MIN FG_CTRL_NUM_MEAS_LOW FG_CTRL_MANY_OUTLIERS FG_CTRL_MARQ FG_CTRL_ROUGHNESS FG_CTRL_FOAM FG_CTRL_ECMWF FG_CTRL_VALID FG_CTRL_NO_SURFACE FG_CTRL_RANGE_ACARD FG_CTRL_SIGMA_ACARD FG_CTRL_USED_FARATEC FG_CTRL_POOR_GEOPHYS FG_CTRL_POOR_RETRIEVAL FG_CTRL_SUSPECT_RFI FG_CTRL_RFI_PRONE_X FG_CTRL_RFI_PRONE_Y FG_CTRL_ADJUSTED_RA FG_CTRL_RETRIEV_FAIL" ;
		string Control_Flags_uncorr:_Unsigned = "true" ;
	ushort Dg_RFI_L1(n_grid_points) ;
		Dg_RFI_L1:_FillValue = 64537US ;
		string Dg_RFI_L1:_Unsigned = "true" ;
	ushort Dg_RFI_X(n_grid_points) ;
		Dg_RFI_X:_FillValue = 64537US ;
		string Dg_RFI_X:_Unsigned = "true" ;
	ushort Dg_RFI_Y(n_grid_points) ;
		Dg_RFI_Y:_FillValue = 64537US ;
		string Dg_RFI_Y:_Unsigned = "true" ;
	ushort Dg_RFI_probability(n_grid_points) ;
		string Dg_RFI_probability:units = "%" ;
		Dg_RFI_probability:_FillValue = 64537US ;
		string Dg_RFI_probability:_Unsigned = "true" ;
	ushort Dg_Suspect_ice(n_grid_points) ;
		Dg_Suspect_ice:_FillValue = 0US ;
		string Dg_Suspect_ice:_Unsigned = "true" ;
	ushort Dg_af_fov(n_grid_points) ;
		Dg_af_fov:_FillValue = 0US ;
		string Dg_af_fov:_Unsigned = "true" ;
	ushort Dg_border_fov(n_grid_points) ;
		Dg_border_fov:_FillValue = 0US ;
		string Dg_border_fov:_Unsigned = "true" ;
	ushort Dg_chi2_Acard(n_grid_points) ;
		Dg_chi2_Acard:_FillValue = 0US ;
		Dg_chi2_Acard:scale_factor = 0.00999999977648258 ;
		Dg_chi2_Acard:scale_offset = 0. ;
		string Dg_chi2_Acard:_Unsigned = "true" ;
	ushort Dg_chi2_P_Acard(n_grid_points) ;
		Dg_chi2_P_Acard:_FillValue = 0US ;
		Dg_chi2_P_Acard:scale_factor = 0.00100000004749745 ;
		Dg_chi2_P_Acard:scale_offset = 0. ;
		string Dg_chi2_P_Acard:_Unsigned = "true" ;
	ushort Dg_chi2_P_corr(n_grid_points) ;
		Dg_chi2_P_corr:_FillValue = 0US ;
		Dg_chi2_P_corr:scale_factor = 0.00100000004749745 ;
		Dg_chi2_P_corr:scale_offset = 0. ;
		string Dg_chi2_P_corr:_Unsigned = "true" ;
	ushort Dg_chi2_P_uncorr(n_grid_points) ;
		Dg_chi2_P_uncorr:_FillValue = 0US ;
		Dg_chi2_P_uncorr:scale_factor = 0.00100000004749745 ;
		Dg_chi2_P_uncorr:scale_offset = 0. ;
		string Dg_chi2_P_uncorr:_Unsigned = "true" ;
	ushort Dg_chi2_corr(n_grid_points) ;
		Dg_chi2_corr:_FillValue = 0US ;
		Dg_chi2_corr:scale_factor = 0.00999999977648258 ;
		Dg_chi2_corr:scale_offset = 0. ;
		string Dg_chi2_corr:_Unsigned = "true" ;
	ushort Dg_chi2_uncorr(n_grid_points) ;
		Dg_chi2_uncorr:_FillValue = 0US ;
		Dg_chi2_uncorr:scale_factor = 0.00999999977648258 ;
		Dg_chi2_uncorr:scale_offset = 0. ;
		string Dg_chi2_uncorr:_Unsigned = "true" ;
	ushort Dg_galactic_Noise_Error(n_grid_points) ;
		Dg_galactic_Noise_Error:_FillValue = 0US ;
		string Dg_galactic_Noise_Error:_Unsigned = "true" ;
	ushort Dg_moonglint(n_grid_points) ;
		Dg_moonglint:_FillValue = 0US ;
		string Dg_moonglint:_Unsigned = "true" ;
	ubyte Dg_num_iter_Acard(n_grid_points) ;
		Dg_num_iter_Acard:_FillValue = 0UB ;
		string Dg_num_iter_Acard:_Unsigned = "true" ;
	ubyte Dg_num_iter_corr(n_grid_points) ;
		Dg_num_iter_corr:_FillValue = 0UB ;
		string Dg_num_iter_corr:_Unsigned = "true" ;
	ubyte Dg_num_iter_uncorr(n_grid_points) ;
		Dg_num_iter_uncorr:_FillValue = 0UB ;
		string Dg_num_iter_uncorr:_Unsigned = "true" ;
	ushort Dg_num_meas_l1c(n_grid_points) ;
		Dg_num_meas_l1c:_FillValue = 0US ;
		string Dg_num_meas_l1c:_Unsigned = "true" ;
	ushort Dg_num_meas_valid(n_grid_points) ;
		Dg_num_meas_valid:_FillValue = 0US ;
		string Dg_num_meas_valid:_Unsigned = "true" ;
	ushort Dg_quality_SSS_anom(n_grid_points) ;
		Dg_quality_SSS_anom:_FillValue = 999US ;
		string Dg_quality_SSS_anom:_Unsigned = "true" ;
	ushort Dg_quality_SSS_corr(n_grid_points) ;
		Dg_quality_SSS_corr:_FillValue = 999US ;
		string Dg_quality_SSS_corr:_Unsigned = "true" ;
	ushort Dg_quality_SSS_uncorr(n_grid_points) ;
		Dg_quality_SSS_uncorr:_FillValue = 999US ;
		string Dg_quality_SSS_uncorr:_Unsigned = "true" ;
	ushort Dg_sky(n_grid_points) ;
		Dg_sky:_FillValue = 64537US ;
		string Dg_sky:_Unsigned = "true" ;
	ushort Dg_sun_glint_L2(n_grid_points) ;
		Dg_sun_glint_L2:_FillValue = 0US ;
		string Dg_sun_glint_L2:_Unsigned = "true" ;
	ushort Dg_sun_glint_area(n_grid_points) ;
		Dg_sun_glint_area:_FillValue = 0US ;
		string Dg_sun_glint_area:_Unsigned = "true" ;
	ushort Dg_sun_glint_fov(n_grid_points) ;
		Dg_sun_glint_fov:_FillValue = 0US ;
		string Dg_sun_glint_fov:_Unsigned = "true" ;
	ushort Dg_sun_tails(n_grid_points) ;
		Dg_sun_tails:_FillValue = 0US ;
		string Dg_sun_tails:_Unsigned = "true" ;
	float Equiv_ftprt_diam(n_grid_points) ;
		string Equiv_ftprt_diam:units = "km" ;
		Equiv_ftprt_diam:_FillValue = -999.f ;
	uint Grid_Point_ID(n_grid_points) ;
		Grid_Point_ID:_FillValue = 0U ;
		string Grid_Point_ID:_Unsigned = "true" ;
	float Latitude(n_grid_points) ;
		string Latitude:units = "deg" ;
		Latitude:_FillValue = -999.f ;
	float Longitude(n_grid_points) ;
		string Longitude:units = "deg" ;
		Longitude:_FillValue = -999.f ;
	float Mean_acq_time(n_grid_points) ;
		string Mean_acq_time:units = "dd" ;
		Mean_acq_time:_FillValue = -999.f ;
	float SSS_anom(n_grid_points) ;
		string SSS_anom:units = "psu" ;
		SSS_anom:_FillValue = -999.f ;
	ushort SSS_climatology(n_grid_points) ;
		SSS_climatology:_FillValue = 0US ;
		SSS_climatology:scale_factor = 0.00999999977648258 ;
		SSS_climatology:scale_offset = 0. ;
		string SSS_climatology:_Unsigned = "true" ;
	float SSS_corr(n_grid_points) ;
		string SSS_corr:units = "psu" ;
		SSS_corr:_FillValue = -999.f ;
	float SSS_uncorr(n_grid_points) ;
		string SSS_uncorr:units = "psu" ;
		SSS_uncorr:_FillValue = -999.f ;
	float SST(n_grid_points) ;
		string SST:units = "°C" ;
		SST:_FillValue = -999.f ;
	uint Science_Flags_Acard(n_grid_points) ;
		Science_Flags_Acard:_FillValue = 0U ;
		Science_Flags_Acard:flag_masks = 1s, 2s, 4s, 8s, 16s, 32s, 64s, 128s, 256s, 512s, 1024s, 2048s, 4096s, 8192s, 16384s, -32768s, 0s, 0s, 0s, 0s, 0s, 0s, 0s ;
		Science_Flags_Acard:flag_values = 1s, 2s, 4s, 8s, 16s, 32s, 64s, 128s, 256s, 512s, 1024s, 2048s, 4096s, 8192s, 16384s, -32768s, 0s, 0s, 0s, 0s, 0s, 0s, 0s ;
		string Science_Flags_Acard:flag_meanings = "FG_SC_LAND_SEA_COAST1 FG_SC_LAND_SEA_COAST2 FG_SC_TEC_GRADIENT FG_SC_IN_CLIM_ICE FG_SC_ICE FG_SC_SUSPECT_ICE FG_SC_RAIN FG_SC_HIGH_WIND FG_SC_LOW_WIND FG_SC_HIGHT_SST FG_SC_LOW_SST FG_SC_HIGH_SSS FG_SC_LOW_SSS FG_SC_SEA_STATE_1 FG_SC_SEA_STATE_2 FG_SC_SEA_STATE_3 FG_SC_SEA_STATE_4 FG_SC_SEA_STATE_5 FG_SC_SEA_STATE_6 FG_SC_SST_FRONT FG_SC_SSS_FRONT FG_SC_ICE_ACARD FG_SC_ECMWF_LAND" ;
		string Science_Flags_Acard:_Unsigned = "true" ;
	uint Science_Flags_anom(n_grid_points) ;
		Science_Flags_anom:_FillValue = 0U ;
		Science_Flags_anom:flag_masks = 1s, 2s, 4s, 8s, 16s, 32s, 64s, 128s, 256s, 512s, 1024s, 2048s, 4096s, 8192s, 16384s, -32768s, 0s, 0s, 0s, 0s, 0s, 0s, 0s ;
		Science_Flags_anom:flag_values = 1s, 2s, 4s, 8s, 16s, 32s, 64s, 128s, 256s, 512s, 1024s, 2048s, 4096s, 8192s, 16384s, -32768s, 0s, 0s, 0s, 0s, 0s, 0s, 0s ;
		string Science_Flags_anom:flag_meanings = "FG_SC_LAND_SEA_COAST1 FG_SC_LAND_SEA_COAST2 FG_SC_TEC_GRADIENT FG_SC_IN_CLIM_ICE FG_SC_ICE FG_SC_SUSPECT_ICE FG_SC_RAIN FG_SC_HIGH_WIND FG_SC_LOW_WIND FG_SC_HIGHT_SST FG_SC_LOW_SST FG_SC_HIGH_SSS FG_SC_LOW_SSS FG_SC_SEA_STATE_1 FG_SC_SEA_STATE_2 FG_SC_SEA_STATE_3 FG_SC_SEA_STATE_4 FG_SC_SEA_STATE_5 FG_SC_SEA_STATE_6 FG_SC_SST_FRONT FG_SC_SSS_FRONT FG_SC_ICE_ACARD FG_SC_ECMWF_LAND" ;
		string Science_Flags_anom:_Unsigned = "true" ;
	uint Science_Flags_corr(n_grid_points) ;
		Science_Flags_corr:_FillValue = 0U ;
		Science_Flags_corr:flag_masks = 1s, 2s, 4s, 8s, 16s, 32s, 64s, 128s, 256s, 512s, 1024s, 2048s, 4096s, 8192s, 16384s, -32768s, 0s, 0s, 0s, 0s, 0s, 0s, 0s ;
		Science_Flags_corr:flag_values = 1s, 2s, 4s, 8s, 16s, 32s, 64s, 128s, 256s, 512s, 1024s, 2048s, 4096s, 8192s, 16384s, -32768s, 0s, 0s, 0s, 0s, 0s, 0s, 0s ;
		string Science_Flags_corr:flag_meanings = "FG_SC_LAND_SEA_COAST1 FG_SC_LAND_SEA_COAST2 FG_SC_TEC_GRADIENT FG_SC_IN_CLIM_ICE FG_SC_ICE FG_SC_SUSPECT_ICE FG_SC_RAIN FG_SC_HIGH_WIND FG_SC_LOW_WIND FG_SC_HIGHT_SST FG_SC_LOW_SST FG_SC_HIGH_SSS FG_SC_LOW_SSS FG_SC_SEA_STATE_1 FG_SC_SEA_STATE_2 FG_SC_SEA_STATE_3 FG_SC_SEA_STATE_4 FG_SC_SEA_STATE_5 FG_SC_SEA_STATE_6 FG_SC_SST_FRONT FG_SC_SSS_FRONT FG_SC_ICE_ACARD FG_SC_ECMWF_LAND" ;
		string Science_Flags_corr:_Unsigned = "true" ;
	uint Science_Flags_uncorr(n_grid_points) ;
		Science_Flags_uncorr:_FillValue = 0U ;
		Science_Flags_uncorr:flag_masks = 1s, 2s, 4s, 8s, 16s, 32s, 64s, 128s, 256s, 512s, 1024s, 2048s, 4096s, 8192s, 16384s, -32768s, 0s, 0s, 0s, 0s, 0s, 0s, 0s ;
		Science_Flags_uncorr:flag_values = 1s, 2s, 4s, 8s, 16s, 32s, 64s, 128s, 256s, 512s, 1024s, 2048s, 4096s, 8192s, 16384s, -32768s, 0s, 0s, 0s, 0s, 0s, 0s, 0s ;
		string Science_Flags_uncorr:flag_meanings = "FG_SC_LAND_SEA_COAST1 FG_SC_LAND_SEA_COAST2 FG_SC_TEC_GRADIENT FG_SC_IN_CLIM_ICE FG_SC_ICE FG_SC_SUSPECT_ICE FG_SC_RAIN FG_SC_HIGH_WIND FG_SC_LOW_WIND FG_SC_HIGHT_SST FG_SC_LOW_SST FG_SC_HIGH_SSS FG_SC_LOW_SSS FG_SC_SEA_STATE_1 FG_SC_SEA_STATE_2 FG_SC_SEA_STATE_3 FG_SC_SEA_STATE_4 FG_SC_SEA_STATE_5 FG_SC_SEA_STATE_6 FG_SC_SST_FRONT FG_SC_SSS_FRONT FG_SC_ICE_ACARD FG_SC_ECMWF_LAND" ;
		string Science_Flags_uncorr:_Unsigned = "true" ;
	float Sigma_Acard(n_grid_points) ;
		Sigma_Acard:_FillValue = -999.f ;
	float Sigma_SSS_anom(n_grid_points) ;
		string Sigma_SSS_anom:units = "psu" ;
		Sigma_SSS_anom:_FillValue = -999.f ;
	float Sigma_SSS_corr(n_grid_points) ;
		string Sigma_SSS_corr:units = "psu" ;
		Sigma_SSS_corr:_FillValue = -999.f ;
	float Sigma_SSS_uncorr(n_grid_points) ;
		string Sigma_SSS_uncorr:units = "psu" ;
		Sigma_SSS_uncorr:_FillValue = -999.f ;
	float Sigma_Tb_42_5H(n_grid_points) ;
		string Sigma_Tb_42_5H:units = "K" ;
		Sigma_Tb_42_5H:_FillValue = -999.f ;
	float Sigma_Tb_42_5V(n_grid_points) ;
		string Sigma_Tb_42_5V:units = "K" ;
		Sigma_Tb_42_5V:_FillValue = -999.f ;
	float Sigma_Tb_42_5X(n_grid_points) ;
		string Sigma_Tb_42_5X:units = "K" ;
		Sigma_Tb_42_5X:_FillValue = -999.f ;
	float Sigma_Tb_42_5Y(n_grid_points) ;
		string Sigma_Tb_42_5Y:units = "K" ;
		Sigma_Tb_42_5Y:_FillValue = -999.f ;
	ushort Sigma_WS_corr(n_grid_points) ;
		Sigma_WS_corr:_FillValue = 0US ;
		Sigma_WS_corr:scale_factor = 0.00100000004749745 ;
		Sigma_WS_corr:scale_offset = 0. ;
		string Sigma_WS_corr:_Unsigned = "true" ;
	float Tb_42_5H(n_grid_points) ;
		string Tb_42_5H:units = "K" ;
		Tb_42_5H:_FillValue = -999.f ;
	float Tb_42_5V(n_grid_points) ;
		string Tb_42_5V:units = "K" ;
		Tb_42_5V:_FillValue = -999.f ;
	float Tb_42_5X(n_grid_points) ;
		string Tb_42_5X:units = "K" ;
		Tb_42_5X:_FillValue = -999.f ;
	float Tb_42_5Y(n_grid_points) ;
		string Tb_42_5Y:units = "K" ;
		Tb_42_5Y:_FillValue = -999.f ;
	float WS(n_grid_points) ;
		string WS:units = "m s-1" ;
		WS:_FillValue = -999.f ;
	ushort WS_corr(n_grid_points) ;
		WS_corr:_FillValue = 0US ;
		WS_corr:scale_factor = 0.00100000004749745 ;
		WS_corr:scale_offset = 0. ;
		string WS_corr:_Unsigned = "true" ;
	float X_swath(n_grid_points) ;
		string X_swath:units = "m" ;
		X_swath:_FillValue = -999.f ;

// global attributes:
		string :creation_date = "UTC=2021-07-01T03:51:46" ;
		string :total_number_of_grid_points = "106350" ;
		string :FH\:File_Name = "SM_OPER_MIR_OSUDP2_20210630T210913_20210630T220228_700_001_1" ;
		string :FH\:File_Description = "L2 Ocean Salinity Output User Data Product." ;
		string :FH\:Notes = "The UDP (User Data Product) is designed for oceanographics and high level centers, it includes geophysical parameters, a theoretical estimate of their accuracy, flags and descriptors of the product quality." ;
		string :FH\:Mission = "SMOS" ;
		string :FH\:File_Class = "OPER" ;
		string :FH\:File_Type = "MIR_OSUDP2" ;
		string :FH\:File_Version = "0001" ;
		string :FH\:Validity_Period\:Validity_Start = "UTC=2021-06-30T21:09:13" ;
		string :FH\:Validity_Period\:Validity_Stop = "UTC=2021-06-30T22:02:28" ;
		string :FH\:Source\:System = "DPGS" ;
		string :FH\:Source\:Creator = "L2OP" ;
		string :FH\:Source\:Creator_Version = "700" ;
		string :FH\:Source\:Creation_Date = "UTC=2021-07-01T03:44:36" ;
		string :VH\:SPH\:QI\:Total_Selected_L1c_Grid_Points = "80650" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:Retrieval_Scheme = "1" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:Land_Rejected = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:Too_Close_To_Land_Rejected = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:Ice_Rejected = "9107" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:Missing_ECMWF_Rejected = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:Too_Few_Measurements_Rejected = "14105" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:Good_Quality_Grid_Points = "49030" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:Poor_Quality_Grid_Points = "10594" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:SQ\:Grid_Point_Type = "Sea" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:SQ\:SSS_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:SQ\:SST_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:SQ\:WS_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:SQ\:Good_Quality = "42416" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:SQ\:Good_Quality_Retrieved = "33881" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:SQ\:Good_Quality_Retrieved_Average_Sigma = "1.300973" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:SQ\:Good_Quality_Failed_Outside_Valid_Range = "138" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:SQ\:Good_Quality_Failed_Sigma_Too_High = "456" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:SQ\:Good_Quality_Failed_Poor_Fit = "7974" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:SQ\:Good_Quality_Failed_Marquardt = "50" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:SQ\:Good_Quality_Failed_Maxiter = "489" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:SQ\:Good_Quality_Failed_OOLUT = "549" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:SQ\:Poor_Quality = "7258" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:SQ\:Poor_Quality_Retrieved = "5481" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:SQ\:Poor_Quality_Retrieved_Average_Sigma = "2.500925" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:NCQ\:Grid_Point_Type = "Near_Coast" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:NCQ\:SSS_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:NCQ\:SST_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:NCQ\:WS_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:NCQ\:Good_Quality = "6614" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:NCQ\:Good_Quality_Retrieved = "3994" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:NCQ\:Good_Quality_Retrieved_Average_Sigma = "2.145041" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:NCQ\:Good_Quality_Failed_Outside_Valid_Range = "331" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:NCQ\:Good_Quality_Failed_Sigma_Too_High = "780" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:NCQ\:Good_Quality_Failed_Poor_Fit = "2270" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:NCQ\:Good_Quality_Failed_Marquardt = "175" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:NCQ\:Good_Quality_Failed_Maxiter = "307" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:NCQ\:Good_Quality_Failed_OOLUT = "993" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:NCQ\:Poor_Quality = "3336" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:NCQ\:Poor_Quality_Retrieved = "2402" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:NCQ\:Poor_Quality_Retrieved_Average_Sigma = "2.491391" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_0\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_0\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_0\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_0\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_0\:Good_Quality = "40" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_0\:Good_Quality_Retrieved = "13" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_0\:Good_Quality_Retrieved_Average_Sigma = "2.271775" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_0\:Good_Quality_Failed_Outside_Valid_Range = "11" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_0\:Good_Quality_Failed_Sigma_Too_High = "13" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_0\:Good_Quality_Failed_Poor_Fit = "26" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_0\:Good_Quality_Failed_Marquardt = "6" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_0\:Good_Quality_Failed_Maxiter = "6" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_0\:Good_Quality_Failed_OOLUT = "14" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_0\:Poor_Quality = "11" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_0\:Poor_Quality_Retrieved = "6" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_0\:Poor_Quality_Retrieved_Average_Sigma = "4.644665" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_1\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_1\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_1\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_1\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_1\:Good_Quality = "32" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_1\:Good_Quality_Retrieved = "25" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_1\:Good_Quality_Retrieved_Average_Sigma = "2.331885" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_1\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_1\:Good_Quality_Failed_Sigma_Too_High = "3" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_1\:Good_Quality_Failed_Poor_Fit = "6" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_1\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_1\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_1\:Good_Quality_Failed_OOLUT = "4" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_1\:Poor_Quality = "185" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_1\:Poor_Quality_Retrieved = "8" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_1\:Poor_Quality_Retrieved_Average_Sigma = "4.768177" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_2\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_2\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_2\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_2\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_2\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_2\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_2\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_2\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_2\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_2\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_2\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_2\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_2\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_2\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_2\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_2\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_3\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_3\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_3\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_3\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_3\:Good_Quality = "6" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_3\:Good_Quality_Retrieved = "6" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_3\:Good_Quality_Retrieved_Average_Sigma = "1.849856" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_3\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_3\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_3\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_3\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_3\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_3\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_3\:Poor_Quality = "92" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_3\:Poor_Quality_Retrieved = "61" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_3\:Poor_Quality_Retrieved_Average_Sigma = "3.938132" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_4\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_4\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_4\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_4\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_4\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_4\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_4\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_4\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_4\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_4\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_4\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_4\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_4\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_4\:Poor_Quality = "371" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_4\:Poor_Quality_Retrieved = "214" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_4\:Poor_Quality_Retrieved_Average_Sigma = "4.211347" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_5\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_5\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_5\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_5\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_5\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_5\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_5\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_5\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_5\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_5\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_5\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_5\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_5\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_5\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_5\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_5\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_6\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_6\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_6\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_6\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_6\:Good_Quality = "127" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_6\:Good_Quality_Retrieved = "36" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_6\:Good_Quality_Retrieved_Average_Sigma = "0.556612" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_6\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_6\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_6\:Good_Quality_Failed_Poor_Fit = "87" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_6\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_6\:Good_Quality_Failed_Maxiter = "9" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_6\:Good_Quality_Failed_OOLUT = "16" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_6\:Poor_Quality = "16" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_6\:Poor_Quality_Retrieved = "9" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_6\:Poor_Quality_Retrieved_Average_Sigma = "3.255918" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_7\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_7\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_7\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_7\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_7\:Good_Quality = "22" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_7\:Good_Quality_Retrieved = "18" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_7\:Good_Quality_Retrieved_Average_Sigma = "0.561522" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_7\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_7\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_7\:Good_Quality_Failed_Poor_Fit = "4" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_7\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_7\:Good_Quality_Failed_Maxiter = "2" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_7\:Good_Quality_Failed_OOLUT = "1" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_7\:Poor_Quality = "17" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_7\:Poor_Quality_Retrieved = "7" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_7\:Poor_Quality_Retrieved_Average_Sigma = "1.677722" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_8\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_8\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_8\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_8\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_8\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_8\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_8\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_8\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_8\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_8\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_8\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_8\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_8\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_8\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_8\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_8\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_9\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_9\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_9\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_9\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_9\:Good_Quality = "273" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_9\:Good_Quality_Retrieved = "160" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_9\:Good_Quality_Retrieved_Average_Sigma = "2.599082" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_9\:Good_Quality_Failed_Outside_Valid_Range = "33" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_9\:Good_Quality_Failed_Sigma_Too_High = "65" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_9\:Good_Quality_Failed_Poor_Fit = "85" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_9\:Good_Quality_Failed_Marquardt = "13" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_9\:Good_Quality_Failed_Maxiter = "32" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_9\:Good_Quality_Failed_OOLUT = "85" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_9\:Poor_Quality = "288" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_9\:Poor_Quality_Retrieved = "240" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_9\:Poor_Quality_Retrieved_Average_Sigma = "3.081223" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_10\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_10\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_10\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_10\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_10\:Good_Quality = "8069" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_10\:Good_Quality_Retrieved = "5269" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_10\:Good_Quality_Retrieved_Average_Sigma = "2.785885" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_10\:Good_Quality_Failed_Outside_Valid_Range = "379" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_10\:Good_Quality_Failed_Sigma_Too_High = "1082" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_10\:Good_Quality_Failed_Poor_Fit = "2346" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_10\:Good_Quality_Failed_Marquardt = "139" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_10\:Good_Quality_Failed_Maxiter = "195" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_10\:Good_Quality_Failed_OOLUT = "1200" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_10\:Poor_Quality = "1600" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_10\:Poor_Quality_Retrieved = "1075" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_10\:Poor_Quality_Retrieved_Average_Sigma = "3.307963" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_11\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_11\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_11\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_11\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_11\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_11\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_11\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_11\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_11\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_11\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_11\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_11\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_11\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_11\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_11\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_11\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_12\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_12\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_12\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_12\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_12\:Good_Quality = "7009" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_12\:Good_Quality_Retrieved = "5885" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_12\:Good_Quality_Retrieved_Average_Sigma = "1.320947" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_12\:Good_Quality_Failed_Outside_Valid_Range = "4" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_12\:Good_Quality_Failed_Sigma_Too_High = "14" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_12\:Good_Quality_Failed_Poor_Fit = "1027" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_12\:Good_Quality_Failed_Marquardt = "48" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_12\:Good_Quality_Failed_Maxiter = "83" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_12\:Good_Quality_Failed_OOLUT = "38" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_12\:Poor_Quality = "1990" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_12\:Poor_Quality_Retrieved = "1563" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_12\:Poor_Quality_Retrieved_Average_Sigma = "2.000069" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_13\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_13\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_13\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_13\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_13\:Good_Quality = "15933" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_13\:Good_Quality_Retrieved = "13481" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_13\:Good_Quality_Retrieved_Average_Sigma = "1.377319" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_13\:Good_Quality_Failed_Outside_Valid_Range = "22" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_13\:Good_Quality_Failed_Sigma_Too_High = "43" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_13\:Good_Quality_Failed_Poor_Fit = "2414" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_13\:Good_Quality_Failed_Marquardt = "5" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_13\:Good_Quality_Failed_Maxiter = "30" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_13\:Good_Quality_Failed_OOLUT = "72" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_13\:Poor_Quality = "3587" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_13\:Poor_Quality_Retrieved = "2944" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_13\:Poor_Quality_Retrieved_Average_Sigma = "2.700215" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_14\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_14\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_14\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_14\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_14\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_14\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_14\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_14\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_14\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_14\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_14\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_14\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_14\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_14\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_14\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_14\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_15\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_15\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_15\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_15\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_15\:Good_Quality = "4315" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_15\:Good_Quality_Retrieved = "2924" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_15\:Good_Quality_Retrieved_Average_Sigma = "0.768287" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_15\:Good_Quality_Failed_Outside_Valid_Range = "18" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_15\:Good_Quality_Failed_Sigma_Too_High = "16" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_15\:Good_Quality_Failed_Poor_Fit = "1107" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_15\:Good_Quality_Failed_Marquardt = "14" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_15\:Good_Quality_Failed_Maxiter = "410" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_15\:Good_Quality_Failed_OOLUT = "52" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_15\:Poor_Quality = "693" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_15\:Poor_Quality_Retrieved = "426" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_15\:Poor_Quality_Retrieved_Average_Sigma = "1.355604" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_16\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_16\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_16\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_16\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_16\:Good_Quality = "13204" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_16\:Good_Quality_Retrieved = "10058" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_16\:Good_Quality_Retrieved_Average_Sigma = "0.878298" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_16\:Good_Quality_Failed_Outside_Valid_Range = "2" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_16\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_16\:Good_Quality_Failed_Poor_Fit = "3142" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_16\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_16\:Good_Quality_Failed_Maxiter = "29" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_16\:Good_Quality_Failed_OOLUT = "60" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_16\:Poor_Quality = "1291" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_16\:Poor_Quality_Retrieved = "989" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_16\:Poor_Quality_Retrieved_Average_Sigma = "1.659203" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_17\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_17\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_17\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_17\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_17\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_17\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_17\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_17\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_17\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_17\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_17\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_17\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_17\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_17\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_17\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_17\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_18\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_18\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_18\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_18\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_18\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_18\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_18\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_18\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_18\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_18\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_18\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_18\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_18\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_18\:Poor_Quality = "12" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_18\:Poor_Quality_Retrieved = "5" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_18\:Poor_Quality_Retrieved_Average_Sigma = "4.724520" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_19\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_19\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_19\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_19\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_19\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_19\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_19\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_19\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_19\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_19\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_19\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_19\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_19\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_19\:Poor_Quality = "7" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_19\:Poor_Quality_Retrieved = "2" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_19\:Poor_Quality_Retrieved_Average_Sigma = "3.689911" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_20\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_20\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_20\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_20\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_20\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_20\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_20\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_20\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_20\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_20\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_20\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_20\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_20\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_20\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_20\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_20\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_21\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_21\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_21\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_21\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_21\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_21\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_21\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_21\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_21\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_21\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_21\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_21\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_21\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_21\:Poor_Quality = "45" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_21\:Poor_Quality_Retrieved = "37" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_21\:Poor_Quality_Retrieved_Average_Sigma = "3.072677" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_22\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_22\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_22\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_22\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_22\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_22\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_22\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_22\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_22\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_22\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_22\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_22\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_22\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_22\:Poor_Quality = "136" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_22\:Poor_Quality_Retrieved = "92" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_22\:Poor_Quality_Retrieved_Average_Sigma = "3.238413" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_23\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_23\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_23\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_23\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_23\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_23\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_23\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_23\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_23\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_23\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_23\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_23\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_23\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_23\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_23\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_23\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_24\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_24\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_24\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_24\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_24\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_24\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_24\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_24\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_24\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_24\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_24\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_24\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_24\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_24\:Poor_Quality = "92" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_24\:Poor_Quality_Retrieved = "72" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_24\:Poor_Quality_Retrieved_Average_Sigma = "1.981403" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_25\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_25\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_25\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_25\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_25\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_25\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_25\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_25\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_25\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_25\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_25\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_25\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_25\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_25\:Poor_Quality = "161" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_25\:Poor_Quality_Retrieved = "133" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_25\:Poor_Quality_Retrieved_Average_Sigma = "2.019211" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_26\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_26\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_26\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_26\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_26\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_26\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_26\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_26\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_26\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_26\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_26\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_26\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_26\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_26\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_26\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_26\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:SIQ\:Grid_Point_Type = "Sea_Ice" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:SIQ\:SSS_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:SIQ\:SST_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:SIQ\:WS_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:SIQ\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:SIQ\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:SIQ\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:SIQ\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:SIQ\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:SIQ\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:SIQ\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:SIQ\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:SIQ\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:SIQ\:Poor_Quality = "41" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:SIQ\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:SIQ\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:Retrieval_Scheme = "2" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:Land_Rejected = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:Too_Close_To_Land_Rejected = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:Ice_Rejected = "9107" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:Missing_ECMWF_Rejected = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:Too_Few_Measurements_Rejected = "14105" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:Good_Quality_Grid_Points = "49030" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:Poor_Quality_Grid_Points = "10594" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:SQ\:Grid_Point_Type = "Sea" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:SQ\:SSS_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:SQ\:SST_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:SQ\:WS_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:SQ\:Good_Quality = "42416" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:SQ\:Good_Quality_Retrieved = "32650" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:SQ\:Good_Quality_Retrieved_Average_Sigma = "1.309669" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:SQ\:Good_Quality_Failed_Outside_Valid_Range = "126" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:SQ\:Good_Quality_Failed_Sigma_Too_High = "467" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:SQ\:Good_Quality_Failed_Poor_Fit = "9129" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:SQ\:Good_Quality_Failed_Marquardt = "66" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:SQ\:Good_Quality_Failed_Maxiter = "638" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:SQ\:Good_Quality_Failed_OOLUT = "573" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:SQ\:Poor_Quality = "7258" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:SQ\:Poor_Quality_Retrieved = "4970" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:SQ\:Poor_Quality_Retrieved_Average_Sigma = "2.602561" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:NCQ\:Grid_Point_Type = "Near_Coast" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:NCQ\:SSS_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:NCQ\:SST_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:NCQ\:WS_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:NCQ\:Good_Quality = "6614" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:NCQ\:Good_Quality_Retrieved = "3196" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:NCQ\:Good_Quality_Retrieved_Average_Sigma = "2.316276" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:NCQ\:Good_Quality_Failed_Outside_Valid_Range = "354" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:NCQ\:Good_Quality_Failed_Sigma_Too_High = "863" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:NCQ\:Good_Quality_Failed_Poor_Fit = "3116" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:NCQ\:Good_Quality_Failed_Marquardt = "226" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:NCQ\:Good_Quality_Failed_Maxiter = "331" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:NCQ\:Good_Quality_Failed_OOLUT = "1302" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:NCQ\:Poor_Quality = "3336" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:NCQ\:Poor_Quality_Retrieved = "2146" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:NCQ\:Poor_Quality_Retrieved_Average_Sigma = "2.596146" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_0\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_0\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_0\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_0\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_0\:Good_Quality = "40" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_0\:Good_Quality_Retrieved = "10" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_0\:Good_Quality_Retrieved_Average_Sigma = "2.410896" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_0\:Good_Quality_Failed_Outside_Valid_Range = "11" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_0\:Good_Quality_Failed_Sigma_Too_High = "13" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_0\:Good_Quality_Failed_Poor_Fit = "29" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_0\:Good_Quality_Failed_Marquardt = "8" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_0\:Good_Quality_Failed_Maxiter = "3" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_0\:Good_Quality_Failed_OOLUT = "17" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_0\:Poor_Quality = "11" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_0\:Poor_Quality_Retrieved = "5" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_0\:Poor_Quality_Retrieved_Average_Sigma = "4.593025" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_1\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_1\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_1\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_1\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_1\:Good_Quality = "32" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_1\:Good_Quality_Retrieved = "23" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_1\:Good_Quality_Retrieved_Average_Sigma = "2.439510" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_1\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_1\:Good_Quality_Failed_Sigma_Too_High = "3" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_1\:Good_Quality_Failed_Poor_Fit = "9" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_1\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_1\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_1\:Good_Quality_Failed_OOLUT = "6" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_1\:Poor_Quality = "185" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_1\:Poor_Quality_Retrieved = "8" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_1\:Poor_Quality_Retrieved_Average_Sigma = "4.803418" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_2\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_2\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_2\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_2\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_2\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_2\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_2\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_2\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_2\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_2\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_2\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_2\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_2\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_2\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_2\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_2\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_3\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_3\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_3\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_3\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_3\:Good_Quality = "6" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_3\:Good_Quality_Retrieved = "6" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_3\:Good_Quality_Retrieved_Average_Sigma = "1.840680" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_3\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_3\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_3\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_3\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_3\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_3\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_3\:Poor_Quality = "92" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_3\:Poor_Quality_Retrieved = "47" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_3\:Poor_Quality_Retrieved_Average_Sigma = "4.075317" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_4\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_4\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_4\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_4\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_4\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_4\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_4\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_4\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_4\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_4\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_4\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_4\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_4\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_4\:Poor_Quality = "371" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_4\:Poor_Quality_Retrieved = "129" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_4\:Poor_Quality_Retrieved_Average_Sigma = "4.287936" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_5\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_5\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_5\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_5\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_5\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_5\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_5\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_5\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_5\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_5\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_5\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_5\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_5\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_5\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_5\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_5\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_6\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_6\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_6\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_6\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_6\:Good_Quality = "127" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_6\:Good_Quality_Retrieved = "28" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_6\:Good_Quality_Retrieved_Average_Sigma = "0.560374" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_6\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_6\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_6\:Good_Quality_Failed_Poor_Fit = "94" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_6\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_6\:Good_Quality_Failed_Maxiter = "28" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_6\:Good_Quality_Failed_OOLUT = "23" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_6\:Poor_Quality = "16" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_6\:Poor_Quality_Retrieved = "1" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_6\:Poor_Quality_Retrieved_Average_Sigma = "1.426370" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_7\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_7\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_7\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_7\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_7\:Good_Quality = "22" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_7\:Good_Quality_Retrieved = "16" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_7\:Good_Quality_Retrieved_Average_Sigma = "0.547665" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_7\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_7\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_7\:Good_Quality_Failed_Poor_Fit = "6" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_7\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_7\:Good_Quality_Failed_Maxiter = "2" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_7\:Good_Quality_Failed_OOLUT = "1" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_7\:Poor_Quality = "17" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_7\:Poor_Quality_Retrieved = "7" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_7\:Poor_Quality_Retrieved_Average_Sigma = "1.832616" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_8\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_8\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_8\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_8\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_8\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_8\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_8\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_8\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_8\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_8\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_8\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_8\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_8\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_8\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_8\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_8\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_9\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_9\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_9\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_9\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_9\:Good_Quality = "273" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_9\:Good_Quality_Retrieved = "155" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_9\:Good_Quality_Retrieved_Average_Sigma = "2.577458" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_9\:Good_Quality_Failed_Outside_Valid_Range = "35" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_9\:Good_Quality_Failed_Sigma_Too_High = "68" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_9\:Good_Quality_Failed_Poor_Fit = "86" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_9\:Good_Quality_Failed_Marquardt = "14" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_9\:Good_Quality_Failed_Maxiter = "34" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_9\:Good_Quality_Failed_OOLUT = "89" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_9\:Poor_Quality = "288" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_9\:Poor_Quality_Retrieved = "244" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_9\:Poor_Quality_Retrieved_Average_Sigma = "3.173979" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_10\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_10\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_10\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_10\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_10\:Good_Quality = "8069" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_10\:Good_Quality_Retrieved = "5009" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_10\:Good_Quality_Retrieved_Average_Sigma = "2.802226" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_10\:Good_Quality_Failed_Outside_Valid_Range = "381" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_10\:Good_Quality_Failed_Sigma_Too_High = "1149" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_10\:Good_Quality_Failed_Poor_Fit = "2608" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_10\:Good_Quality_Failed_Marquardt = "146" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_10\:Good_Quality_Failed_Maxiter = "192" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_10\:Good_Quality_Failed_OOLUT = "1331" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_10\:Poor_Quality = "1600" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_10\:Poor_Quality_Retrieved = "1041" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_10\:Poor_Quality_Retrieved_Average_Sigma = "3.312484" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_11\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_11\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_11\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_11\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_11\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_11\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_11\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_11\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_11\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_11\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_11\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_11\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_11\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_11\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_11\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_11\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_12\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_12\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_12\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_12\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_12\:Good_Quality = "7009" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_12\:Good_Quality_Retrieved = "5553" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_12\:Good_Quality_Retrieved_Average_Sigma = "1.349544" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_12\:Good_Quality_Failed_Outside_Valid_Range = "8" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_12\:Good_Quality_Failed_Sigma_Too_High = "19" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_12\:Good_Quality_Failed_Poor_Fit = "1358" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_12\:Good_Quality_Failed_Marquardt = "70" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_12\:Good_Quality_Failed_Maxiter = "126" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_12\:Good_Quality_Failed_OOLUT = "68" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_12\:Poor_Quality = "1990" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_12\:Poor_Quality_Retrieved = "1438" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_12\:Poor_Quality_Retrieved_Average_Sigma = "2.169792" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_13\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_13\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_13\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_13\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_13\:Good_Quality = "15933" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_13\:Good_Quality_Retrieved = "12618" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_13\:Good_Quality_Retrieved_Average_Sigma = "1.389448" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_13\:Good_Quality_Failed_Outside_Valid_Range = "16" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_13\:Good_Quality_Failed_Sigma_Too_High = "48" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_13\:Good_Quality_Failed_Poor_Fit = "3254" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_13\:Good_Quality_Failed_Marquardt = "11" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_13\:Good_Quality_Failed_Maxiter = "79" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_13\:Good_Quality_Failed_OOLUT = "214" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_13\:Poor_Quality = "3587" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_13\:Poor_Quality_Retrieved = "2533" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_13\:Poor_Quality_Retrieved_Average_Sigma = "2.911479" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_14\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_14\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_14\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_14\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_14\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_14\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_14\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_14\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_14\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_14\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_14\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_14\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_14\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_14\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_14\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_14\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_15\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_15\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_15\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_15\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_15\:Good_Quality = "4315" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_15\:Good_Quality_Retrieved = "2837" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_15\:Good_Quality_Retrieved_Average_Sigma = "0.767496" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_15\:Good_Quality_Failed_Outside_Valid_Range = "29" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_15\:Good_Quality_Failed_Sigma_Too_High = "30" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_15\:Good_Quality_Failed_Poor_Fit = "1196" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_15\:Good_Quality_Failed_Marquardt = "43" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_15\:Good_Quality_Failed_Maxiter = "474" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_15\:Good_Quality_Failed_OOLUT = "67" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_15\:Poor_Quality = "693" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_15\:Poor_Quality_Retrieved = "404" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_15\:Poor_Quality_Retrieved_Average_Sigma = "1.257553" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_16\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_16\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_16\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_16\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_16\:Good_Quality = "13204" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_16\:Good_Quality_Retrieved = "9591" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_16\:Good_Quality_Retrieved_Average_Sigma = "0.876707" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_16\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_16\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_16\:Good_Quality_Failed_Poor_Fit = "3605" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_16\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_16\:Good_Quality_Failed_Maxiter = "31" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_16\:Good_Quality_Failed_OOLUT = "59" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_16\:Poor_Quality = "1291" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_16\:Poor_Quality_Retrieved = "907" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_16\:Poor_Quality_Retrieved_Average_Sigma = "1.710565" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_17\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_17\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_17\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_17\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_17\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_17\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_17\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_17\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_17\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_17\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_17\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_17\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_17\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_17\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_17\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_17\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_18\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_18\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_18\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_18\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_18\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_18\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_18\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_18\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_18\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_18\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_18\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_18\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_18\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_18\:Poor_Quality = "12" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_18\:Poor_Quality_Retrieved = "5" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_18\:Poor_Quality_Retrieved_Average_Sigma = "4.715192" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_19\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_19\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_19\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_19\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_19\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_19\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_19\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_19\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_19\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_19\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_19\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_19\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_19\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_19\:Poor_Quality = "7" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_19\:Poor_Quality_Retrieved = "2" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_19\:Poor_Quality_Retrieved_Average_Sigma = "3.695637" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_20\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_20\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_20\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_20\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_20\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_20\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_20\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_20\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_20\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_20\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_20\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_20\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_20\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_20\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_20\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_20\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_21\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_21\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_21\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_21\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_21\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_21\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_21\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_21\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_21\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_21\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_21\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_21\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_21\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_21\:Poor_Quality = "45" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_21\:Poor_Quality_Retrieved = "34" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_21\:Poor_Quality_Retrieved_Average_Sigma = "3.077266" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_22\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_22\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_22\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_22\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_22\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_22\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_22\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_22\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_22\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_22\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_22\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_22\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_22\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_22\:Poor_Quality = "136" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_22\:Poor_Quality_Retrieved = "104" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_22\:Poor_Quality_Retrieved_Average_Sigma = "3.421102" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_23\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_23\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_23\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_23\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_23\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_23\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_23\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_23\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_23\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_23\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_23\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_23\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_23\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_23\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_23\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_23\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_24\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_24\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_24\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_24\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_24\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_24\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_24\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_24\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_24\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_24\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_24\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_24\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_24\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_24\:Poor_Quality = "92" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_24\:Poor_Quality_Retrieved = "74" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_24\:Poor_Quality_Retrieved_Average_Sigma = "2.013027" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_25\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_25\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_25\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_25\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_25\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_25\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_25\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_25\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_25\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_25\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_25\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_25\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_25\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_25\:Poor_Quality = "161" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_25\:Poor_Quality_Retrieved = "133" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_25\:Poor_Quality_Retrieved_Average_Sigma = "2.016223" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_26\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_26\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_26\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_26\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_26\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_26\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_26\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_26\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_26\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_26\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_26\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_26\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_26\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_26\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_26\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_26\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:SIQ\:Grid_Point_Type = "Sea_Ice" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:SIQ\:SSS_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:SIQ\:SST_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:SIQ\:WS_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:SIQ\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:SIQ\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:SIQ\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:SIQ\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:SIQ\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:SIQ\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:SIQ\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:SIQ\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:SIQ\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:SIQ\:Poor_Quality = "41" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:SIQ\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:SIQ\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:Retrieval_Scheme = "3" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:Land_Rejected = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:Too_Close_To_Land_Rejected = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:Ice_Rejected = "9107" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:Missing_ECMWF_Rejected = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:Too_Few_Measurements_Rejected = "14105" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:Good_Quality_Grid_Points = "49030" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:Poor_Quality_Grid_Points = "10594" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:SQ\:Grid_Point_Type = "Sea" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:SQ\:SSS_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:SQ\:SST_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:SQ\:WS_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:SQ\:Good_Quality = "42416" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:SQ\:Good_Quality_Retrieved = "33881" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:SQ\:Good_Quality_Retrieved_Average_Sigma = "1.300973" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:SQ\:Good_Quality_Failed_Outside_Valid_Range = "138" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:SQ\:Good_Quality_Failed_Sigma_Too_High = "456" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:SQ\:Good_Quality_Failed_Poor_Fit = "7974" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:SQ\:Good_Quality_Failed_Marquardt = "50" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:SQ\:Good_Quality_Failed_Maxiter = "489" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:SQ\:Good_Quality_Failed_OOLUT = "549" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:SQ\:Poor_Quality = "7258" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:SQ\:Poor_Quality_Retrieved = "5481" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:SQ\:Poor_Quality_Retrieved_Average_Sigma = "2.500925" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:NCQ\:Grid_Point_Type = "Near_Coast" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:NCQ\:SSS_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:NCQ\:SST_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:NCQ\:WS_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:NCQ\:Good_Quality = "6614" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:NCQ\:Good_Quality_Retrieved = "3994" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:NCQ\:Good_Quality_Retrieved_Average_Sigma = "2.145041" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:NCQ\:Good_Quality_Failed_Outside_Valid_Range = "331" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:NCQ\:Good_Quality_Failed_Sigma_Too_High = "780" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:NCQ\:Good_Quality_Failed_Poor_Fit = "2270" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:NCQ\:Good_Quality_Failed_Marquardt = "175" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:NCQ\:Good_Quality_Failed_Maxiter = "307" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:NCQ\:Good_Quality_Failed_OOLUT = "993" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:NCQ\:Poor_Quality = "3336" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:NCQ\:Poor_Quality_Retrieved = "2402" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:NCQ\:Poor_Quality_Retrieved_Average_Sigma = "2.491391" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_0\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_0\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_0\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_0\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_0\:Good_Quality = "40" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_0\:Good_Quality_Retrieved = "13" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_0\:Good_Quality_Retrieved_Average_Sigma = "2.271775" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_0\:Good_Quality_Failed_Outside_Valid_Range = "11" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_0\:Good_Quality_Failed_Sigma_Too_High = "13" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_0\:Good_Quality_Failed_Poor_Fit = "26" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_0\:Good_Quality_Failed_Marquardt = "6" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_0\:Good_Quality_Failed_Maxiter = "6" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_0\:Good_Quality_Failed_OOLUT = "14" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_0\:Poor_Quality = "11" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_0\:Poor_Quality_Retrieved = "6" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_0\:Poor_Quality_Retrieved_Average_Sigma = "4.644665" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_1\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_1\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_1\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_1\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_1\:Good_Quality = "32" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_1\:Good_Quality_Retrieved = "25" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_1\:Good_Quality_Retrieved_Average_Sigma = "2.331885" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_1\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_1\:Good_Quality_Failed_Sigma_Too_High = "3" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_1\:Good_Quality_Failed_Poor_Fit = "6" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_1\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_1\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_1\:Good_Quality_Failed_OOLUT = "4" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_1\:Poor_Quality = "185" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_1\:Poor_Quality_Retrieved = "8" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_1\:Poor_Quality_Retrieved_Average_Sigma = "4.768177" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_2\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_2\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_2\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_2\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_2\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_2\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_2\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_2\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_2\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_2\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_2\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_2\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_2\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_2\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_2\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_2\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_3\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_3\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_3\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_3\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_3\:Good_Quality = "6" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_3\:Good_Quality_Retrieved = "6" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_3\:Good_Quality_Retrieved_Average_Sigma = "1.849856" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_3\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_3\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_3\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_3\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_3\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_3\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_3\:Poor_Quality = "92" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_3\:Poor_Quality_Retrieved = "61" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_3\:Poor_Quality_Retrieved_Average_Sigma = "3.938132" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_4\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_4\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_4\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_4\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_4\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_4\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_4\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_4\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_4\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_4\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_4\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_4\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_4\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_4\:Poor_Quality = "371" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_4\:Poor_Quality_Retrieved = "214" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_4\:Poor_Quality_Retrieved_Average_Sigma = "4.211347" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_5\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_5\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_5\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_5\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_5\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_5\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_5\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_5\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_5\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_5\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_5\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_5\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_5\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_5\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_5\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_5\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_6\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_6\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_6\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_6\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_6\:Good_Quality = "127" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_6\:Good_Quality_Retrieved = "36" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_6\:Good_Quality_Retrieved_Average_Sigma = "0.556612" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_6\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_6\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_6\:Good_Quality_Failed_Poor_Fit = "87" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_6\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_6\:Good_Quality_Failed_Maxiter = "9" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_6\:Good_Quality_Failed_OOLUT = "16" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_6\:Poor_Quality = "16" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_6\:Poor_Quality_Retrieved = "9" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_6\:Poor_Quality_Retrieved_Average_Sigma = "3.255918" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_7\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_7\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_7\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_7\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_7\:Good_Quality = "22" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_7\:Good_Quality_Retrieved = "18" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_7\:Good_Quality_Retrieved_Average_Sigma = "0.561522" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_7\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_7\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_7\:Good_Quality_Failed_Poor_Fit = "4" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_7\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_7\:Good_Quality_Failed_Maxiter = "2" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_7\:Good_Quality_Failed_OOLUT = "1" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_7\:Poor_Quality = "17" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_7\:Poor_Quality_Retrieved = "7" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_7\:Poor_Quality_Retrieved_Average_Sigma = "1.677722" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_8\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_8\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_8\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_8\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_8\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_8\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_8\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_8\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_8\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_8\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_8\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_8\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_8\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_8\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_8\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_8\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_9\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_9\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_9\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_9\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_9\:Good_Quality = "273" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_9\:Good_Quality_Retrieved = "160" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_9\:Good_Quality_Retrieved_Average_Sigma = "2.599082" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_9\:Good_Quality_Failed_Outside_Valid_Range = "33" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_9\:Good_Quality_Failed_Sigma_Too_High = "65" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_9\:Good_Quality_Failed_Poor_Fit = "85" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_9\:Good_Quality_Failed_Marquardt = "13" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_9\:Good_Quality_Failed_Maxiter = "32" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_9\:Good_Quality_Failed_OOLUT = "85" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_9\:Poor_Quality = "288" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_9\:Poor_Quality_Retrieved = "240" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_9\:Poor_Quality_Retrieved_Average_Sigma = "3.081223" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_10\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_10\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_10\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_10\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_10\:Good_Quality = "8069" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_10\:Good_Quality_Retrieved = "5269" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_10\:Good_Quality_Retrieved_Average_Sigma = "2.785885" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_10\:Good_Quality_Failed_Outside_Valid_Range = "379" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_10\:Good_Quality_Failed_Sigma_Too_High = "1082" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_10\:Good_Quality_Failed_Poor_Fit = "2346" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_10\:Good_Quality_Failed_Marquardt = "139" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_10\:Good_Quality_Failed_Maxiter = "195" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_10\:Good_Quality_Failed_OOLUT = "1200" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_10\:Poor_Quality = "1600" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_10\:Poor_Quality_Retrieved = "1075" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_10\:Poor_Quality_Retrieved_Average_Sigma = "3.307963" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_11\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_11\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_11\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_11\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_11\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_11\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_11\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_11\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_11\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_11\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_11\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_11\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_11\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_11\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_11\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_11\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_12\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_12\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_12\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_12\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_12\:Good_Quality = "7009" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_12\:Good_Quality_Retrieved = "5885" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_12\:Good_Quality_Retrieved_Average_Sigma = "1.320947" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_12\:Good_Quality_Failed_Outside_Valid_Range = "4" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_12\:Good_Quality_Failed_Sigma_Too_High = "14" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_12\:Good_Quality_Failed_Poor_Fit = "1027" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_12\:Good_Quality_Failed_Marquardt = "48" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_12\:Good_Quality_Failed_Maxiter = "83" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_12\:Good_Quality_Failed_OOLUT = "38" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_12\:Poor_Quality = "1990" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_12\:Poor_Quality_Retrieved = "1563" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_12\:Poor_Quality_Retrieved_Average_Sigma = "2.000069" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_13\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_13\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_13\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_13\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_13\:Good_Quality = "15933" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_13\:Good_Quality_Retrieved = "13481" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_13\:Good_Quality_Retrieved_Average_Sigma = "1.377319" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_13\:Good_Quality_Failed_Outside_Valid_Range = "22" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_13\:Good_Quality_Failed_Sigma_Too_High = "43" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_13\:Good_Quality_Failed_Poor_Fit = "2414" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_13\:Good_Quality_Failed_Marquardt = "5" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_13\:Good_Quality_Failed_Maxiter = "30" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_13\:Good_Quality_Failed_OOLUT = "72" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_13\:Poor_Quality = "3587" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_13\:Poor_Quality_Retrieved = "2944" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_13\:Poor_Quality_Retrieved_Average_Sigma = "2.700215" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_14\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_14\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_14\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_14\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_14\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_14\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_14\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_14\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_14\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_14\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_14\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_14\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_14\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_14\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_14\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_14\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_15\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_15\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_15\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_15\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_15\:Good_Quality = "4315" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_15\:Good_Quality_Retrieved = "2924" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_15\:Good_Quality_Retrieved_Average_Sigma = "0.768287" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_15\:Good_Quality_Failed_Outside_Valid_Range = "18" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_15\:Good_Quality_Failed_Sigma_Too_High = "16" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_15\:Good_Quality_Failed_Poor_Fit = "1107" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_15\:Good_Quality_Failed_Marquardt = "14" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_15\:Good_Quality_Failed_Maxiter = "410" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_15\:Good_Quality_Failed_OOLUT = "52" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_15\:Poor_Quality = "693" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_15\:Poor_Quality_Retrieved = "426" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_15\:Poor_Quality_Retrieved_Average_Sigma = "1.355604" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_16\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_16\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_16\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_16\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_16\:Good_Quality = "13204" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_16\:Good_Quality_Retrieved = "10058" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_16\:Good_Quality_Retrieved_Average_Sigma = "0.878298" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_16\:Good_Quality_Failed_Outside_Valid_Range = "2" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_16\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_16\:Good_Quality_Failed_Poor_Fit = "3142" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_16\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_16\:Good_Quality_Failed_Maxiter = "29" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_16\:Good_Quality_Failed_OOLUT = "60" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_16\:Poor_Quality = "1291" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_16\:Poor_Quality_Retrieved = "989" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_16\:Poor_Quality_Retrieved_Average_Sigma = "1.659203" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_17\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_17\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_17\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_17\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_17\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_17\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_17\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_17\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_17\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_17\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_17\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_17\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_17\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_17\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_17\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_17\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_18\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_18\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_18\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_18\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_18\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_18\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_18\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_18\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_18\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_18\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_18\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_18\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_18\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_18\:Poor_Quality = "12" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_18\:Poor_Quality_Retrieved = "5" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_18\:Poor_Quality_Retrieved_Average_Sigma = "4.724520" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_19\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_19\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_19\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_19\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_19\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_19\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_19\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_19\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_19\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_19\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_19\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_19\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_19\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_19\:Poor_Quality = "7" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_19\:Poor_Quality_Retrieved = "2" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_19\:Poor_Quality_Retrieved_Average_Sigma = "3.689911" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_20\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_20\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_20\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_20\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_20\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_20\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_20\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_20\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_20\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_20\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_20\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_20\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_20\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_20\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_20\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_20\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_21\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_21\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_21\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_21\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_21\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_21\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_21\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_21\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_21\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_21\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_21\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_21\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_21\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_21\:Poor_Quality = "45" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_21\:Poor_Quality_Retrieved = "37" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_21\:Poor_Quality_Retrieved_Average_Sigma = "3.072677" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_22\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_22\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_22\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_22\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_22\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_22\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_22\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_22\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_22\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_22\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_22\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_22\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_22\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_22\:Poor_Quality = "136" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_22\:Poor_Quality_Retrieved = "92" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_22\:Poor_Quality_Retrieved_Average_Sigma = "3.238413" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_23\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_23\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_23\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_23\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_23\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_23\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_23\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_23\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_23\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_23\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_23\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_23\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_23\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_23\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_23\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_23\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_24\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_24\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_24\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_24\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_24\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_24\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_24\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_24\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_24\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_24\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_24\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_24\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_24\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_24\:Poor_Quality = "92" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_24\:Poor_Quality_Retrieved = "72" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_24\:Poor_Quality_Retrieved_Average_Sigma = "1.981403" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_25\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_25\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_25\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_25\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_25\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_25\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_25\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_25\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_25\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_25\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_25\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_25\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_25\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_25\:Poor_Quality = "161" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_25\:Poor_Quality_Retrieved = "133" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_25\:Poor_Quality_Retrieved_Average_Sigma = "2.019211" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_26\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_26\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_26\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_26\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_26\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_26\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_26\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_26\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_26\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_26\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_26\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_26\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_26\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_26\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_26\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_26\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:SIQ\:Grid_Point_Type = "Sea_Ice" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:SIQ\:SSS_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:SIQ\:SST_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:SIQ\:WS_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:SIQ\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:SIQ\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:SIQ\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:SIQ\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:SIQ\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:SIQ\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:SIQ\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:SIQ\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:SIQ\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:SIQ\:Poor_Quality = "41" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:SIQ\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:SIQ\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:Retrieval_Scheme = "4" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:Land_Rejected = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:Too_Close_To_Land_Rejected = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:Ice_Rejected = "9107" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:Missing_ECMWF_Rejected = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:Too_Few_Measurements_Rejected = "14105" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:Good_Quality_Grid_Points = "49030" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:Poor_Quality_Grid_Points = "10594" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:SQ\:Grid_Point_Type = "Sea" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:SQ\:SSS_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:SQ\:SST_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:SQ\:WS_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:SQ\:Good_Quality = "42416" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:SQ\:Good_Quality_Retrieved = "38092" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:SQ\:Good_Quality_Retrieved_Average_Sigma = "0.777640" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:SQ\:Good_Quality_Failed_Outside_Valid_Range = "725" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:SQ\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:SQ\:Good_Quality_Failed_Poor_Fit = "3680" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:SQ\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:SQ\:Good_Quality_Failed_Maxiter = "5" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:SQ\:Good_Quality_Failed_OOLUT = "3670" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:SQ\:Poor_Quality = "7258" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:SQ\:Poor_Quality_Retrieved = "5930" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:SQ\:Poor_Quality_Retrieved_Average_Sigma = "1.312244" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:NCQ\:Grid_Point_Type = "Near_Coast" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:NCQ\:SSS_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:NCQ\:SST_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:NCQ\:WS_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:NCQ\:Good_Quality = "6614" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:NCQ\:Good_Quality_Retrieved = "5275" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:NCQ\:Good_Quality_Retrieved_Average_Sigma = "0.713190" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:NCQ\:Good_Quality_Failed_Outside_Valid_Range = "108" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:NCQ\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:NCQ\:Good_Quality_Failed_Poor_Fit = "1336" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:NCQ\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:NCQ\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:NCQ\:Good_Quality_Failed_OOLUT = "1330" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:NCQ\:Poor_Quality = "3336" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:NCQ\:Poor_Quality_Retrieved = "2822" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:NCQ\:Poor_Quality_Retrieved_Average_Sigma = "1.012104" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_0\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_0\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_0\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_0\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_0\:Good_Quality = "40" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_0\:Good_Quality_Retrieved = "31" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_0\:Good_Quality_Retrieved_Average_Sigma = "0.584082" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_0\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_0\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_0\:Good_Quality_Failed_Poor_Fit = "9" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_0\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_0\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_0\:Good_Quality_Failed_OOLUT = "9" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_0\:Poor_Quality = "11" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_0\:Poor_Quality_Retrieved = "11" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_0\:Poor_Quality_Retrieved_Average_Sigma = "1.497783" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_1\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_1\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_1\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_1\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_1\:Good_Quality = "32" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_1\:Good_Quality_Retrieved = "30" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_1\:Good_Quality_Retrieved_Average_Sigma = "0.623371" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_1\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_1\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_1\:Good_Quality_Failed_Poor_Fit = "2" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_1\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_1\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_1\:Good_Quality_Failed_OOLUT = "2" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_1\:Poor_Quality = "185" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_1\:Poor_Quality_Retrieved = "120" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_1\:Poor_Quality_Retrieved_Average_Sigma = "1.599651" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_2\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_2\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_2\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_2\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_2\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_2\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_2\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_2\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_2\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_2\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_2\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_2\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_2\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_2\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_2\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_2\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_3\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_3\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_3\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_3\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_3\:Good_Quality = "6" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_3\:Good_Quality_Retrieved = "6" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_3\:Good_Quality_Retrieved_Average_Sigma = "0.953346" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_3\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_3\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_3\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_3\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_3\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_3\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_3\:Poor_Quality = "92" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_3\:Poor_Quality_Retrieved = "72" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_3\:Poor_Quality_Retrieved_Average_Sigma = "1.688501" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_4\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_4\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_4\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_4\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_4\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_4\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_4\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_4\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_4\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_4\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_4\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_4\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_4\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_4\:Poor_Quality = "371" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_4\:Poor_Quality_Retrieved = "314" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_4\:Poor_Quality_Retrieved_Average_Sigma = "1.663750" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_5\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_5\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_5\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_5\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_5\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_5\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_5\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_5\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_5\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_5\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_5\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_5\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_5\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_5\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_5\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_5\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_6\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_6\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_6\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_6\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_6\:Good_Quality = "127" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_6\:Good_Quality_Retrieved = "48" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_6\:Good_Quality_Retrieved_Average_Sigma = "0.726662" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_6\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_6\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_6\:Good_Quality_Failed_Poor_Fit = "79" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_6\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_6\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_6\:Good_Quality_Failed_OOLUT = "79" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_6\:Poor_Quality = "16" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_6\:Poor_Quality_Retrieved = "9" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_6\:Poor_Quality_Retrieved_Average_Sigma = "1.440257" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_7\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_7\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_7\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_7\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_7\:Good_Quality = "22" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_7\:Good_Quality_Retrieved = "18" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_7\:Good_Quality_Retrieved_Average_Sigma = "0.760549" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_7\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_7\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_7\:Good_Quality_Failed_Poor_Fit = "4" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_7\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_7\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_7\:Good_Quality_Failed_OOLUT = "4" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_7\:Poor_Quality = "17" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_7\:Poor_Quality_Retrieved = "6" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_7\:Poor_Quality_Retrieved_Average_Sigma = "1.655105" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_8\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_8\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_8\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_8\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_8\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_8\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_8\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_8\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_8\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_8\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_8\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_8\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_8\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_8\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_8\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_8\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_9\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_9\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_9\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_9\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_9\:Good_Quality = "273" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_9\:Good_Quality_Retrieved = "228" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_9\:Good_Quality_Retrieved_Average_Sigma = "0.667519" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_9\:Good_Quality_Failed_Outside_Valid_Range = "1" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_9\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_9\:Good_Quality_Failed_Poor_Fit = "44" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_9\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_9\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_9\:Good_Quality_Failed_OOLUT = "45" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_9\:Poor_Quality = "288" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_9\:Poor_Quality_Retrieved = "249" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_9\:Poor_Quality_Retrieved_Average_Sigma = "1.094154" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_10\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_10\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_10\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_10\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_10\:Good_Quality = "8069" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_10\:Good_Quality_Retrieved = "6840" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_10\:Good_Quality_Retrieved_Average_Sigma = "0.689680" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_10\:Good_Quality_Failed_Outside_Valid_Range = "83" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_10\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_10\:Good_Quality_Failed_Poor_Fit = "1224" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_10\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_10\:Good_Quality_Failed_Maxiter = "5" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_10\:Good_Quality_Failed_OOLUT = "1229" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_10\:Poor_Quality = "1600" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_10\:Poor_Quality_Retrieved = "1347" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_10\:Poor_Quality_Retrieved_Average_Sigma = "1.023891" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_11\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_11\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_11\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_11\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_11\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_11\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_11\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_11\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_11\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_11\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_11\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_11\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_11\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_11\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_11\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_11\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_12\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_12\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_12\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_12\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_12\:Good_Quality = "7009" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_12\:Good_Quality_Retrieved = "6588" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_12\:Good_Quality_Retrieved_Average_Sigma = "0.757073" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_12\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_12\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_12\:Good_Quality_Failed_Poor_Fit = "421" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_12\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_12\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_12\:Good_Quality_Failed_OOLUT = "414" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_12\:Poor_Quality = "1990" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_12\:Poor_Quality_Retrieved = "1804" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_12\:Poor_Quality_Retrieved_Average_Sigma = "0.902115" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_13\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_13\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_13\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_13\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_13\:Good_Quality = "15933" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_13\:Good_Quality_Retrieved = "14872" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_13\:Good_Quality_Retrieved_Average_Sigma = "0.744029" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_13\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_13\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_13\:Good_Quality_Failed_Poor_Fit = "1061" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_13\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_13\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_13\:Good_Quality_Failed_OOLUT = "1017" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_13\:Poor_Quality = "3587" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_13\:Poor_Quality_Retrieved = "3124" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_13\:Poor_Quality_Retrieved_Average_Sigma = "1.219597" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_14\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_14\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_14\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_14\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_14\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_14\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_14\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_14\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_14\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_14\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_14\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_14\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_14\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_14\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_14\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_14\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_15\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_15\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_15\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_15\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_15\:Good_Quality = "4315" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_15\:Good_Quality_Retrieved = "3022" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_15\:Good_Quality_Retrieved_Average_Sigma = "0.822249" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_15\:Good_Quality_Failed_Outside_Valid_Range = "694" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_15\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_15\:Good_Quality_Failed_Poor_Fit = "675" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_15\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_15\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_15\:Good_Quality_Failed_OOLUT = "1096" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_15\:Poor_Quality = "693" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_15\:Poor_Quality_Retrieved = "418" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_15\:Poor_Quality_Retrieved_Average_Sigma = "1.274173" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_16\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_16\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_16\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_16\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_16\:Good_Quality = "13204" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_16\:Good_Quality_Retrieved = "11684" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_16\:Good_Quality_Retrieved_Average_Sigma = "0.846080" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_16\:Good_Quality_Failed_Outside_Valid_Range = "55" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_16\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_16\:Good_Quality_Failed_Poor_Fit = "1497" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_16\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_16\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_16\:Good_Quality_Failed_OOLUT = "1105" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_16\:Poor_Quality = "1291" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_16\:Poor_Quality_Retrieved = "996" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_16\:Poor_Quality_Retrieved_Average_Sigma = "1.601620" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_17\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_17\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_17\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_17\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_17\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_17\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_17\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_17\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_17\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_17\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_17\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_17\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_17\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_17\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_17\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_17\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_18\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_18\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_18\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_18\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_18\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_18\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_18\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_18\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_18\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_18\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_18\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_18\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_18\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_18\:Poor_Quality = "12" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_18\:Poor_Quality_Retrieved = "9" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_18\:Poor_Quality_Retrieved_Average_Sigma = "1.653254" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_19\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_19\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_19\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_19\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_19\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_19\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_19\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_19\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_19\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_19\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_19\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_19\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_19\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_19\:Poor_Quality = "7" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_19\:Poor_Quality_Retrieved = "6" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_19\:Poor_Quality_Retrieved_Average_Sigma = "1.644945" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_20\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_20\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_20\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_20\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_20\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_20\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_20\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_20\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_20\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_20\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_20\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_20\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_20\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_20\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_20\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_20\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_21\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_21\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_21\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_21\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_21\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_21\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_21\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_21\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_21\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_21\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_21\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_21\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_21\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_21\:Poor_Quality = "45" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_21\:Poor_Quality_Retrieved = "41" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_21\:Poor_Quality_Retrieved_Average_Sigma = "1.816824" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_22\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_22\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_22\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_22\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_22\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_22\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_22\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_22\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_22\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_22\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_22\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_22\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_22\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_22\:Poor_Quality = "136" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_22\:Poor_Quality_Retrieved = "102" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_22\:Poor_Quality_Retrieved_Average_Sigma = "1.893596" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_23\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_23\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_23\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_23\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_23\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_23\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_23\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_23\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_23\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_23\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_23\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_23\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_23\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_23\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_23\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_23\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_24\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_24\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_24\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_24\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_24\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_24\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_24\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_24\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_24\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_24\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_24\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_24\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_24\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_24\:Poor_Quality = "92" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_24\:Poor_Quality_Retrieved = "31" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_24\:Poor_Quality_Retrieved_Average_Sigma = "2.030431" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_25\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_25\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_25\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_25\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_25\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_25\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_25\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_25\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_25\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_25\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_25\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_25\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_25\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_25\:Poor_Quality = "161" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_25\:Poor_Quality_Retrieved = "93" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_25\:Poor_Quality_Retrieved_Average_Sigma = "2.045601" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_26\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_26\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_26\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_26\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_26\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_26\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_26\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_26\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_26\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_26\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_26\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_26\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_26\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_26\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_26\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_26\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:SIQ\:Grid_Point_Type = "Sea_Ice" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:SIQ\:SSS_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:SIQ\:SST_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:SIQ\:WS_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:SIQ\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:SIQ\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:SIQ\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:SIQ\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:SIQ\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:SIQ\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:SIQ\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:SIQ\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:SIQ\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:SIQ\:Poor_Quality = "41" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:SIQ\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:SIQ\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_0\:Retrieved_Parameter_0\:name = "SSS" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_0\:Retrieved_Parameter_0\:unit = "Practical Salinity Unit (PSU)" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_0\:Retrieved_Parameter_0\:description = "Surface salinity of the sea at gridpoint" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_0\:Retrieved_Parameter_1\:name = "SST" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_0\:Retrieved_Parameter_1\:unit = "Kelvin" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_0\:Retrieved_Parameter_1\:description = "Surface temperature of the sea at gridpoint" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_0\:Retrieved_Parameter_2\:name = "UN10" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_0\:Retrieved_Parameter_2\:unit = "m.s-1" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_0\:Retrieved_Parameter_2\:description = "U component of neutral wind 10m above surface" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_0\:Retrieved_Parameter_3\:name = "VN10" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_0\:Retrieved_Parameter_3\:unit = "m.s-1" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_0\:Retrieved_Parameter_3\:description = "V component of neutral wind 10m above surface" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_0\:Retrieved_Parameter_4\:name = "tec" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_0\:Retrieved_Parameter_4\:unit = "tecu" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_0\:Retrieved_Parameter_4\:description = "Total Electronic Content of the ionosphere below SMOS" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_0\:Retrieved_Parameter_5\:name = "not used" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_0\:Retrieved_Parameter_5\:unit = "none" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_0\:Retrieved_Parameter_5\:description = "no parameter defined" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_0\:Retrieved_Parameter_6\:name = "not used" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_0\:Retrieved_Parameter_6\:unit = "none" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_0\:Retrieved_Parameter_6\:description = "no parameter defined" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_0\:Retrieved_Parameter_7\:name = "not used" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_0\:Retrieved_Parameter_7\:unit = "none" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_0\:Retrieved_Parameter_7\:description = "no parameter defined" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_0\:Retrieved_Parameter_8\:name = "not used" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_0\:Retrieved_Parameter_8\:unit = "none" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_0\:Retrieved_Parameter_8\:description = "no parameter defined" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_0\:Retrieved_Parameter_9\:name = "not used" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_0\:Retrieved_Parameter_9\:unit = "none" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_0\:Retrieved_Parameter_9\:description = "no parameter defined" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_1\:Retrieved_Parameter_0\:name = "SSS" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_1\:Retrieved_Parameter_0\:unit = "Practical Salinity Unit (PSU)" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_1\:Retrieved_Parameter_0\:description = "Surface salinity of the sea at gridpoint" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_1\:Retrieved_Parameter_1\:name = "SST" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_1\:Retrieved_Parameter_1\:unit = "Kelvin" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_1\:Retrieved_Parameter_1\:description = "Surface temperature of the sea at gridpoint" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_1\:Retrieved_Parameter_2\:name = "UN10" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_1\:Retrieved_Parameter_2\:unit = "m.s-1" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_1\:Retrieved_Parameter_2\:description = "U component of neutral wind 10m above surface" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_1\:Retrieved_Parameter_3\:name = "VN10" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_1\:Retrieved_Parameter_3\:unit = "m.s-1" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_1\:Retrieved_Parameter_3\:description = "V component of neutral wind 10m above surface" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_1\:Retrieved_Parameter_4\:name = "tec" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_1\:Retrieved_Parameter_4\:unit = "tecu" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_1\:Retrieved_Parameter_4\:description = "Total Electronic Content of the ionosphere below SMOS" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_1\:Retrieved_Parameter_5\:name = "not used" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_1\:Retrieved_Parameter_5\:unit = "none" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_1\:Retrieved_Parameter_5\:description = "no parameter defined" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_1\:Retrieved_Parameter_6\:name = "not used" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_1\:Retrieved_Parameter_6\:unit = "none" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_1\:Retrieved_Parameter_6\:description = "no parameter defined" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_1\:Retrieved_Parameter_7\:name = "not used" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_1\:Retrieved_Parameter_7\:unit = "none" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_1\:Retrieved_Parameter_7\:description = "no parameter defined" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_1\:Retrieved_Parameter_8\:name = "not used" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_1\:Retrieved_Parameter_8\:unit = "none" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_1\:Retrieved_Parameter_8\:description = "no parameter defined" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_1\:Retrieved_Parameter_9\:name = "not used" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_1\:Retrieved_Parameter_9\:unit = "none" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_1\:Retrieved_Parameter_9\:description = "no parameter defined" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_2\:Retrieved_Parameter_0\:name = "SSS" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_2\:Retrieved_Parameter_0\:unit = "Practical Salinity Unit (PSU)" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_2\:Retrieved_Parameter_0\:description = "Surface salinity of the sea at gridpoint" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_2\:Retrieved_Parameter_1\:name = "SST" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_2\:Retrieved_Parameter_1\:unit = "Kelvin" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_2\:Retrieved_Parameter_1\:description = "Surface temperature of the sea at gridpoint" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_2\:Retrieved_Parameter_2\:name = "UN10" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_2\:Retrieved_Parameter_2\:unit = "m.s-1" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_2\:Retrieved_Parameter_2\:description = "U component of neutral wind 10m above surface" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_2\:Retrieved_Parameter_3\:name = "VN10" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_2\:Retrieved_Parameter_3\:unit = "m.s-1" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_2\:Retrieved_Parameter_3\:description = "V component of neutral wind 10m above surface" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_2\:Retrieved_Parameter_4\:name = "tec" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_2\:Retrieved_Parameter_4\:unit = "tecu" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_2\:Retrieved_Parameter_4\:description = "Total Electronic Content of the ionosphere below SMOS" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_2\:Retrieved_Parameter_5\:name = "not used" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_2\:Retrieved_Parameter_5\:unit = "none" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_2\:Retrieved_Parameter_5\:description = "no parameter defined" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_2\:Retrieved_Parameter_6\:name = "not used" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_2\:Retrieved_Parameter_6\:unit = "none" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_2\:Retrieved_Parameter_6\:description = "no parameter defined" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_2\:Retrieved_Parameter_7\:name = "not used" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_2\:Retrieved_Parameter_7\:unit = "none" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_2\:Retrieved_Parameter_7\:description = "no parameter defined" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_2\:Retrieved_Parameter_8\:name = "not used" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_2\:Retrieved_Parameter_8\:unit = "none" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_2\:Retrieved_Parameter_8\:description = "no parameter defined" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_2\:Retrieved_Parameter_9\:name = "not used" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_2\:Retrieved_Parameter_9\:unit = "none" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_2\:Retrieved_Parameter_9\:description = "no parameter defined" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_3\:Retrieved_Parameter_0\:name = "Acard" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_3\:Retrieved_Parameter_0\:unit = "dl" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_3\:Retrieved_Parameter_0\:description = "Acard coefficient for cardioid model" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_3\:Retrieved_Parameter_1\:name = "SST" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_3\:Retrieved_Parameter_1\:unit = "Kelvin" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_3\:Retrieved_Parameter_1\:description = "Surface temperature of the sea at gridpoint" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_3\:Retrieved_Parameter_2\:name = "not used" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_3\:Retrieved_Parameter_2\:unit = "none" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_3\:Retrieved_Parameter_2\:description = "no parameter defined" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_3\:Retrieved_Parameter_3\:name = "not used" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_3\:Retrieved_Parameter_3\:unit = "none" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_3\:Retrieved_Parameter_3\:description = "no parameter defined" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_3\:Retrieved_Parameter_4\:name = "not used" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_3\:Retrieved_Parameter_4\:unit = "none" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_3\:Retrieved_Parameter_4\:description = "no parameter defined" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_3\:Retrieved_Parameter_5\:name = "not used" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_3\:Retrieved_Parameter_5\:unit = "none" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_3\:Retrieved_Parameter_5\:description = "no parameter defined" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_3\:Retrieved_Parameter_6\:name = "not used" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_3\:Retrieved_Parameter_6\:unit = "none" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_3\:Retrieved_Parameter_6\:description = "no parameter defined" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_3\:Retrieved_Parameter_7\:name = "not used" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_3\:Retrieved_Parameter_7\:unit = "none" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_3\:Retrieved_Parameter_7\:description = "no parameter defined" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_3\:Retrieved_Parameter_8\:name = "not used" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_3\:Retrieved_Parameter_8\:unit = "none" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_3\:Retrieved_Parameter_8\:description = "no parameter defined" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_3\:Retrieved_Parameter_9\:name = "not used" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_3\:Retrieved_Parameter_9\:unit = "none" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_3\:Retrieved_Parameter_9\:description = "no parameter defined" ;
		string :VH\:SPH\:MI\:SPH_Descriptor = "MIR_OSUDP2_SPH" ;
		string :VH\:SPH\:MI\:Checksum = "2323233818" ;
		string :VH\:SPH\:MI\:Header_Schema = "HDR_SM_XXXX_MIR_OSUDP2_0400.xsd" ;
		string :VH\:SPH\:MI\:Datablock_Schema = "DBL_SM_XXXX_MIR_OSUDP2_0401.binXschema.xml" ;
		string :VH\:SPH\:MI\:Header_Size = "168709" ;
		string :VH\:SPH\:MI\:Datablock_Size = "00020206504" ;
		string :VH\:SPH\:MI\:HW_Identifier = "0003" ;
		string :VH\:SPH\:MI\:TI\:Precise_Validity_Start = "UTC=2021-06-30T21:09:12.434579" ;
		string :VH\:SPH\:MI\:TI\:Precise_Validity_Stop = "UTC=2021-06-30T22:02:28.074411" ;
		string :VH\:SPH\:MI\:TI\:Abs_Orbit_Start = "+61281" ;
		string :VH\:SPH\:MI\:TI\:Start_Time_ANX_T = "1286.293116" ;
		string :VH\:SPH\:MI\:TI\:Abs_Orbit_Stop = "+61281" ;
		string :VH\:SPH\:MI\:TI\:Stop_Time_ANX_T = "4481.932948" ;
		string :VH\:SPH\:MI\:TI\:UTC_at_ANX = "UTC=2021-06-30T20:47:46.141463" ;
		string :VH\:SPH\:MI\:TI\:Long_at_ANX = "+138.381497" ;
		string :VH\:SPH\:MI\:TI\:Ascending_Flag = "D" ;
		string :VH\:SPH\:MI\:TI\:Polarisation_Flag = "F" ;
		string :VH\:SPH\:LODS\:Data_Set_0\:DS_Name = "SSS_SWATH" ;
		string :VH\:SPH\:LODS\:Data_Set_0\:DS_Type = "M" ;
		string :VH\:SPH\:LODS\:Data_Set_0\:DS_Size = "0020206504" ;
		string :VH\:SPH\:LODS\:Data_Set_0\:DS_Offset = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_0\:Num_DSR = "0000106350" ;
		string :VH\:SPH\:LODS\:Data_Set_0\:DSR_Size = "00000190" ;
		string :VH\:SPH\:LODS\:Data_Set_0\:Byte_Order = "0123" ;
		string :VH\:SPH\:LODS\:Data_Set_1\:DS_Name = "L1C_OS_FILE" ;
		string :VH\:SPH\:LODS\:Data_Set_1\:DS_Type = "R" ;
		string :VH\:SPH\:LODS\:Data_Set_1\:DS_Size = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_1\:DS_Offset = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_1\:Ref_Filename = "SM_OPER_MIR_SCSF1C_20210630T210913_20210630T220228_724_001_1" ;
		string :VH\:SPH\:LODS\:Data_Set_1\:Num_DSR = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_1\:DSR_Size = "00000000" ;
		string :VH\:SPH\:LODS\:Data_Set_1\:Byte_Order = "0000" ;
		string :VH\:SPH\:LODS\:Data_Set_2\:DS_Name = "DGG_FILE" ;
		string :VH\:SPH\:LODS\:Data_Set_2\:DS_Type = "R" ;
		string :VH\:SPH\:LODS\:Data_Set_2\:DS_Size = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_2\:DS_Offset = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_2\:Ref_Filename = "SM_OPER_AUX_DGG____20050101T000000_20500101T000000_300_003_3" ;
		string :VH\:SPH\:LODS\:Data_Set_2\:Num_DSR = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_2\:DSR_Size = "00000000" ;
		string :VH\:SPH\:LODS\:Data_Set_2\:Byte_Order = "0000" ;
		string :VH\:SPH\:LODS\:Data_Set_3\:DS_Name = "IERS_BULLETIN_B_FILE" ;
		string :VH\:SPH\:LODS\:Data_Set_3\:DS_Type = "R" ;
		string :VH\:SPH\:LODS\:Data_Set_3\:DS_Size = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_3\:DS_Offset = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_3\:Ref_Filename = "SM_OPER_AUX_BULL_B_20210402T000000_20500101T000000_120_001_3" ;
		string :VH\:SPH\:LODS\:Data_Set_3\:Num_DSR = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_3\:DSR_Size = "00000000" ;
		string :VH\:SPH\:LODS\:Data_Set_3\:Byte_Order = "0000" ;
		string :VH\:SPH\:LODS\:Data_Set_4\:DS_Name = "BESTFITPLANE_FILE" ;
		string :VH\:SPH\:LODS\:Data_Set_4\:DS_Type = "R" ;
		string :VH\:SPH\:LODS\:Data_Set_4\:DS_Size = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_4\:DS_Offset = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_4\:Ref_Filename = "SM_OPER_AUX_BFP____20050101T000000_20500101T000000_340_004_3" ;
		string :VH\:SPH\:LODS\:Data_Set_4\:Num_DSR = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_4\:DSR_Size = "00000000" ;
		string :VH\:SPH\:LODS\:Data_Set_4\:Byte_Order = "0000" ;
		string :VH\:SPH\:LODS\:Data_Set_5\:DS_Name = "MISPOINTING_FILE" ;
		string :VH\:SPH\:LODS\:Data_Set_5\:DS_Type = "R" ;
		string :VH\:SPH\:LODS\:Data_Set_5\:DS_Size = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_5\:DS_Offset = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_5\:Ref_Filename = "SM_OPER_AUX_MISP___20050101T000000_20500101T000000_300_004_3" ;
		string :VH\:SPH\:LODS\:Data_Set_5\:Num_DSR = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_5\:DSR_Size = "00000000" ;
		string :VH\:SPH\:LODS\:Data_Set_5\:Byte_Order = "0000" ;
		string :VH\:SPH\:LODS\:Data_Set_6\:DS_Name = "ECMWF_FILE" ;
		string :VH\:SPH\:LODS\:Data_Set_6\:DS_Type = "R" ;
		string :VH\:SPH\:LODS\:Data_Set_6\:DS_Size = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_6\:DS_Offset = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_6\:Ref_Filename = "SM_OPER_AUX_ECMWF__20210630T210900_20210630T221540_318_001_3" ;
		string :VH\:SPH\:LODS\:Data_Set_6\:Num_DSR = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_6\:DSR_Size = "00000000" ;
		string :VH\:SPH\:LODS\:Data_Set_6\:Byte_Order = "0000" ;
		string :VH\:SPH\:LODS\:Data_Set_7\:DS_Name = "FLAT_SEA_FILE" ;
		string :VH\:SPH\:LODS\:Data_Set_7\:DS_Type = "R" ;
		string :VH\:SPH\:LODS\:Data_Set_7\:DS_Size = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_7\:DS_Offset = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_7\:Ref_Filename = "SM_OPER_AUX_FLTSEA_20050101T000000_20500101T000000_001_012_3" ;
		string :VH\:SPH\:LODS\:Data_Set_7\:Num_DSR = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_7\:DSR_Size = "00000000" ;
		string :VH\:SPH\:LODS\:Data_Set_7\:Byte_Order = "0000" ;
		string :VH\:SPH\:LODS\:Data_Set_8\:DS_Name = "ROUGHNESS_IPSL_FILE" ;
		string :VH\:SPH\:LODS\:Data_Set_8\:DS_Type = "R" ;
		string :VH\:SPH\:LODS\:Data_Set_8\:DS_Size = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_8\:DS_Offset = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_8\:Ref_Filename = "SM_OPER_AUX_RGHNS1_20050101T000000_20500101T000000_001_016_3" ;
		string :VH\:SPH\:LODS\:Data_Set_8\:Num_DSR = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_8\:DSR_Size = "00000000" ;
		string :VH\:SPH\:LODS\:Data_Set_8\:Byte_Order = "0000" ;
		string :VH\:SPH\:LODS\:Data_Set_9\:DS_Name = "ROUGHNESS_IFREMER_FILE" ;
		string :VH\:SPH\:LODS\:Data_Set_9\:DS_Type = "R" ;
		string :VH\:SPH\:LODS\:Data_Set_9\:DS_Size = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_9\:DS_Offset = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_9\:Ref_Filename = "SM_OPER_AUX_RGHNS2_20050101T000000_20500101T000000_001_013_3" ;
		string :VH\:SPH\:LODS\:Data_Set_9\:Num_DSR = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_9\:DSR_Size = "00000000" ;
		string :VH\:SPH\:LODS\:Data_Set_9\:Byte_Order = "0000" ;
		string :VH\:SPH\:LODS\:Data_Set_10\:DS_Name = "ROUGHNESS_ICM_CSIC_FILE" ;
		string :VH\:SPH\:LODS\:Data_Set_10\:DS_Type = "R" ;
		string :VH\:SPH\:LODS\:Data_Set_10\:DS_Size = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_10\:DS_Offset = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_10\:Ref_Filename = "SM_OPER_AUX_RGHNS3_20050101T000000_20500101T000000_001_016_3" ;
		string :VH\:SPH\:LODS\:Data_Set_10\:Num_DSR = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_10\:DSR_Size = "00000000" ;
		string :VH\:SPH\:LODS\:Data_Set_10\:Byte_Order = "0000" ;
		string :VH\:SPH\:LODS\:Data_Set_11\:DS_Name = "GALAXY_OS_FILE" ;
		string :VH\:SPH\:LODS\:Data_Set_11\:DS_Type = "R" ;
		string :VH\:SPH\:LODS\:Data_Set_11\:DS_Size = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_11\:DS_Offset = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_11\:Ref_Filename = "SM_OPER_AUX_GAL_OS_20050101T000000_20500101T000000_001_011_3" ;
		string :VH\:SPH\:LODS\:Data_Set_11\:Num_DSR = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_11\:DSR_Size = "00000000" ;
		string :VH\:SPH\:LODS\:Data_Set_11\:Byte_Order = "0000" ;
		string :VH\:SPH\:LODS\:Data_Set_12\:DS_Name = "GALAXY_2OS_FILE" ;
		string :VH\:SPH\:LODS\:Data_Set_12\:DS_Type = "R" ;
		string :VH\:SPH\:LODS\:Data_Set_12\:DS_Size = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_12\:DS_Offset = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_12\:Ref_Filename = "SM_OPER_AUX_GAL2OS_20050101T000000_20500101T000000_001_016_3" ;
		string :VH\:SPH\:LODS\:Data_Set_12\:Num_DSR = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_12\:DSR_Size = "00000000" ;
		string :VH\:SPH\:LODS\:Data_Set_12\:Byte_Order = "0000" ;
		string :VH\:SPH\:LODS\:Data_Set_13\:DS_Name = "SUNGLINT_FILE" ;
		string :VH\:SPH\:LODS\:Data_Set_13\:DS_Type = "R" ;
		string :VH\:SPH\:LODS\:Data_Set_13\:DS_Size = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_13\:DS_Offset = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_13\:Ref_Filename = "SM_OPER_AUX_SGLINT_20050101T000000_20500101T000000_001_012_3" ;
		string :VH\:SPH\:LODS\:Data_Set_13\:Num_DSR = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_13\:DSR_Size = "00000000" ;
		string :VH\:SPH\:LODS\:Data_Set_13\:Byte_Order = "0000" ;
		string :VH\:SPH\:LODS\:Data_Set_14\:DS_Name = "ATMOS_FILE" ;
		string :VH\:SPH\:LODS\:Data_Set_14\:DS_Type = "R" ;
		string :VH\:SPH\:LODS\:Data_Set_14\:DS_Size = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_14\:DS_Offset = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_14\:Ref_Filename = "SM_OPER_AUX_ATMOS__20050101T000000_20500101T000000_001_010_3" ;
		string :VH\:SPH\:LODS\:Data_Set_14\:Num_DSR = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_14\:DSR_Size = "00000000" ;
		string :VH\:SPH\:LODS\:Data_Set_14\:Byte_Order = "0000" ;
		string :VH\:SPH\:LODS\:Data_Set_15\:DS_Name = "DISTAN_FILE" ;
		string :VH\:SPH\:LODS\:Data_Set_15\:DS_Type = "R" ;
		string :VH\:SPH\:LODS\:Data_Set_15\:DS_Size = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_15\:DS_Offset = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_15\:Ref_Filename = "SM_OPER_AUX_DISTAN_20050101T000000_20500101T000000_001_011_3" ;
		string :VH\:SPH\:LODS\:Data_Set_15\:Num_DSR = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_15\:DSR_Size = "00000000" ;
		string :VH\:SPH\:LODS\:Data_Set_15\:Byte_Order = "0000" ;
		string :VH\:SPH\:LODS\:Data_Set_16\:DS_Name = "CLIMATOLOGY_SSS_FILE" ;
		string :VH\:SPH\:LODS\:Data_Set_16\:DS_Type = "R" ;
		string :VH\:SPH\:LODS\:Data_Set_16\:DS_Size = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_16\:DS_Offset = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_16\:Ref_Filename = "SM_OPER_AUX_SSS____20050101T000000_20500101T000000_001_014_3" ;
		string :VH\:SPH\:LODS\:Data_Set_16\:Num_DSR = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_16\:DSR_Size = "00000000" ;
		string :VH\:SPH\:LODS\:Data_Set_16\:Byte_Order = "0000" ;
		string :VH\:SPH\:LODS\:Data_Set_17\:DS_Name = "CLIMATOLOGY_SSSCLI_FILE" ;
		string :VH\:SPH\:LODS\:Data_Set_17\:DS_Type = "R" ;
		string :VH\:SPH\:LODS\:Data_Set_17\:DS_Size = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_17\:DS_Offset = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_17\:Ref_Filename = "SM_OPER_AUX_SSSCLI_20050101T000000_20500101T000000_001_002_3" ;
		string :VH\:SPH\:LODS\:Data_Set_17\:Num_DSR = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_17\:DSR_Size = "00000000" ;
		string :VH\:SPH\:LODS\:Data_Set_17\:Byte_Order = "0000" ;
		string :VH\:SPH\:LODS\:Data_Set_18\:DS_Name = "OCEAN_SALINITY_CONFIG_FILE" ;
		string :VH\:SPH\:LODS\:Data_Set_18\:DS_Type = "R" ;
		string :VH\:SPH\:LODS\:Data_Set_18\:DS_Size = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_18\:DS_Offset = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_18\:Ref_Filename = "SM_OPER_AUX_CNFOSF_20050101T000000_20500101T000000_001_032_3" ;
		string :VH\:SPH\:LODS\:Data_Set_18\:Num_DSR = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_18\:DSR_Size = "00000000" ;
		string :VH\:SPH\:LODS\:Data_Set_18\:Byte_Order = "0000" ;
		string :VH\:SPH\:LODS\:Data_Set_19\:DS_Name = "OTT1F_FILE" ;
		string :VH\:SPH\:LODS\:Data_Set_19\:DS_Type = "R" ;
		string :VH\:SPH\:LODS\:Data_Set_19\:DS_Size = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_19\:DS_Offset = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_19\:Ref_Filename = "SM_OPER_AUX_OTT1F__20210624T082406_20500101T000000_700_001_1" ;
		string :VH\:SPH\:LODS\:Data_Set_19\:Num_DSR = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_19\:DSR_Size = "00000000" ;
		string :VH\:SPH\:LODS\:Data_Set_19\:Byte_Order = "0000" ;
		string :VH\:SPH\:LODS\:Data_Set_20\:DS_Name = "OTT2F_FILE" ;
		string :VH\:SPH\:LODS\:Data_Set_20\:DS_Type = "R" ;
		string :VH\:SPH\:LODS\:Data_Set_20\:DS_Size = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_20\:DS_Offset = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_20\:Ref_Filename = "SM_OPER_AUX_OTT2F__20210624T082406_20500101T000000_700_001_1" ;
		string :VH\:SPH\:LODS\:Data_Set_20\:Num_DSR = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_20\:DSR_Size = "00000000" ;
		string :VH\:SPH\:LODS\:Data_Set_20\:Byte_Order = "0000" ;
		string :VH\:SPH\:LODS\:Data_Set_21\:DS_Name = "OTT3F_FILE" ;
		string :VH\:SPH\:LODS\:Data_Set_21\:DS_Type = "R" ;
		string :VH\:SPH\:LODS\:Data_Set_21\:DS_Size = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_21\:DS_Offset = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_21\:Ref_Filename = "SM_OPER_AUX_OTT3F__20210624T082406_20500101T000000_700_001_1" ;
		string :VH\:SPH\:LODS\:Data_Set_21\:Num_DSR = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_21\:DSR_Size = "00000000" ;
		string :VH\:SPH\:LODS\:Data_Set_21\:Byte_Order = "0000" ;
		string :VH\:SPH\:LODS\:Data_Set_22\:DS_Name = "DGGRFI_FILE" ;
		string :VH\:SPH\:LODS\:Data_Set_22\:DS_Type = "R" ;
		string :VH\:SPH\:LODS\:Data_Set_22\:DS_Size = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_22\:DS_Offset = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_22\:Ref_Filename = "SM_OPER_AUX_DGGRFI_20210629T000711_20500101T000000_600_001_1" ;
		string :VH\:SPH\:LODS\:Data_Set_22\:Num_DSR = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_22\:DSR_Size = "00000000" ;
		string :VH\:SPH\:LODS\:Data_Set_22\:Byte_Order = "0000" ;
		string :VH\:SPH\:LODS\:Data_Set_23\:DS_Name = "MIXED_SCENE_OTT_FILE" ;
		string :VH\:SPH\:LODS\:Data_Set_23\:DS_Type = "R" ;
		string :VH\:SPH\:LODS\:Data_Set_23\:DS_Size = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_23\:DS_Offset = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_23\:Ref_Filename = "SM_OPER_AUX_MSOTT__20050101T000000_20500101T000000_001_002_3" ;
		string :VH\:SPH\:LODS\:Data_Set_23\:Num_DSR = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_23\:DSR_Size = "00000000" ;
		string :VH\:SPH\:LODS\:Data_Set_23\:Byte_Order = "0000" ;
		string :VH\:SPH\:L2PL\:Start_Lat = "+075.719335" ;
		string :VH\:SPH\:L2PL\:Start_Long = "+097.548779" ;
		string :VH\:SPH\:L2PL\:Stop_Lat = "-081.598965" ;
		string :VH\:SPH\:L2PL\:Stop_Long = "-150.028234" ;
		string :VH\:SPH\:L2PL\:Mid_Lat = "+005.419643" ;
		string :VH\:SPH\:L2PL\:Mid_Lon = "-052.859901" ;
		string :VH\:SPH\:L2PL\:Southernmost_Latitude = "-067.069000" ;
		string :VH\:SPH\:L2PL\:Southernmost_Gridpoint_ID = "6166549" ;
		string :VH\:SPH\:L2PL\:Northernmost_Latitude = "+079.646004" ;
		string :VH\:SPH\:L2PL\:Northernmost_Gridpoint_ID = "0002902" ;
		string :VH\:SPH\:L2PL\:Easternmost_Longitude = "+049.222000" ;
		string :VH\:SPH\:L2PL\:Easternmost_Gridpoint_ID = "4084941" ;
		string :VH\:SPH\:L2PL\:Westernmost_Longitude = "-090.652000" ;
		string :VH\:SPH\:L2PL\:Westernmost_Gridpoint_ID = "6155252" ;
		string :VH\:MPH\:Ref_Doc = "SO-TN-IDR-GS-0006" ;
		string :VH\:MPH\:Acquisition_Station = "SVLD" ;
		string :VH\:MPH\:Processing_Centre = "ESAC" ;
		string :VH\:MPH\:Logical_Proc_Centre = "FPC" ;
		string :VH\:MPH\:Product_Confidence = "NOMINAL" ;
		string :VH\:MPH\:OI\:Phase = "+001" ;
		string :VH\:MPH\:OI\:Cycle = "+037" ;
		string :VH\:MPH\:OI\:Rel_Orbit = "+01161" ;
		string :VH\:MPH\:OI\:Abs_Orbit = "+61281" ;
		string :VH\:MPH\:OI\:OSV_TAI = "TAI=2021-06-30T21:08:37.000000" ;
		string :VH\:MPH\:OI\:OSV_UTC = "UTC=2021-06-30T21:08:00.000000" ;
		string :VH\:MPH\:OI\:OSV_UT1 = "UT1=2021-06-30T21:08:00.590000" ;
		string :VH\:MPH\:OI\:X_Position = "-0616039.695" ;
		string :VH\:MPH\:OI\:Y_Position = "+2121521.304" ;
		string :VH\:MPH\:OI\:Z_Position = "+6778739.127" ;
		string :VH\:MPH\:OI\:X_Velocity = "+5304.621980" ;
		string :VH\:MPH\:OI\:Y_Velocity = "-4977.113140" ;
		string :VH\:MPH\:OI\:Z_Velocity = "+2035.575410" ;
		string :VH\:MPH\:OI\:Vector_Source = "FP" ;
		:history = "Mon Sep 25 18:31:09 2023: ncks -d n_grid_points,100,100000,2000 /scratch1/NCEPDEV/stmp4/Shastri.Paturi/forAndrew/gdas.20210701/00/SSS/SM_OPER_MIR_OSUDP2_20210630T210913_20210630T220228_700_001_1.nc sss_smos_1" ;
		:NCO = "netCDF Operators version 5.0.6 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco)" ;
data:

 A_card = _, _, _, _, 47.31788, _, _, _, 46.17867, 51.31869, 49.9962, _, 
    50.43442, 50.62265, _, _, 55.63542, 57.76852, 50.0545, _, 62.13977, 
    58.59171, 60.83137, _, 63.83729, 62.17725, 63.68936, 61.53354, 62.58694, 
    59.6455, 59.03718, 62.53212, _, 62.65478, _, _, _, _, 51.13051, 51.49137, 
    50.58967, _, _, 49.71899, 48.04662, 48.08532, 48.52538, _, _, _ ;

 Coast_distance = 21, 10, 4, 8, 12, _, _, _, 4, 25, 4, _, 30, 45, 13, 60, 39, 
    41, 13, 24, 61, 42, 47, 48, 85, 83, 62, 44, 47, 41, 32, 56, 49, 24, _, _, 
    _, 8, 7, 22, 11, _, _, 16, 8, 29, 27, 19, 1, _ ;

 Control_Flags_Acard = 437420040, 437420040, 437420040, 437420040, 411468288, 
    50468865, 453115905, 50468865, 143032832, 411468288, 411468288, 50468865, 
    411468288, 8815104, 453122049, 453122048, 8815104, 8815104, 428249600, 
    50468865, 411468288, 8815104, 8815104, 453122048, 411467776, 411468288, 
    411468288, 445022728, 411468288, 445022984, 411468288, 42369544, 
    50468864, 428249600, 50468865, 50468865, 50468865, 184686593, 8815104, 
    428249856, 411468544, 50462721, 50468865, 8815104, 159814144, 8815104, 
    25596416, 402817536, 184680449, 184680449 ;

 Control_Flags_anom = 453148672, 453148672, 453148672, 453148672, 445023792, 
    50468865, 453115905, 50468865, 176587312, 445023776, 411468320, 50468865, 
    411468320, 8815104, 453122049, 453155328, 8815104, 8815104, 428249632, 
    50468865, 411468288, 8815104, 8815104, 453155328, 411467776, 411468288, 
    411468288, 445022744, 411468288, 445023032, 411468288, 42369592, 
    50502144, 495358496, 50468865, 50468865, 50468865, 184686593, 8815136, 
    428249888, 411468576, 50462721, 50468865, 8815136, 159814176, 8815136, 
    25596416, 453149184, 184680449, 251789313 ;

 Control_Flags_corr = 453148672, 453148672, 453148672, 453148672, 445023792, 
    50468865, 453115905, 50468865, 176587312, 445023776, 411468320, 50468865, 
    411468320, 8815104, 453122049, 453155328, 8815104, 8815104, 428249632, 
    50468865, 411468288, 8815104, 8815104, 453155328, 411467776, 411468288, 
    411468288, 445022744, 411468288, 445023032, 411468288, 42369592, 
    50502144, 495358496, 50468865, 50468865, 50468865, 184686593, 8815136, 
    428249888, 411468576, 50462721, 50468865, 8815136, 159814176, 8815136, 
    25596416, 453149184, 184680449, 251789313 ;

 Control_Flags_uncorr = 453115904, 453115904, 453115904, 453115904, 
    445023280, 50468865, 453115905, 50468865, 176586800, 411467808, 
    411467808, 50468865, 411467808, 8814592, 453122049, 453122048, 8814592, 
    8814592, 428249120, 50468865, 411467776, 8814592, 8814592, 453122048, 
    411467776, 411467776, 411467776, 445022232, 445022224, 445022520, 
    411467776, 42369080, 50468864, 495357984, 50468865, 50468865, 50468865, 
    184686593, 42369072, 428249376, 411468064, 50462721, 50468865, 8814624, 
    159813664, 8814624, 25595904, 453115904, 184680449, 251789313 ;

 Dg_RFI_L1 = 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0 ;

 Dg_RFI_X = 2, 13, 4, 0, 13, 0, 15, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 0, 0, 0, 0, 3, 3, 0, 0, 0, 0, 0, 
    0, 0, 29, 0, 64 ;

 Dg_RFI_Y = 1, 11, 2, 0, 14, 0, 18, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 0, 0, 0, 0, 3, 2, 0, 0, 0, 0, 0, 
    0, 0, 26, 0, 65 ;

 Dg_RFI_probability = 24, 37, 4, 3, 42, 0, 4, 0, 2, 8, 3, 0, 2, 2, 3, 13, 1, 
    1, 3, 2, 3, 2, 2, 2, 5, 4, 3, 4, 4, 2, 7, 1, 2, 8, 0, 0, 0, 2, 1, 3, 2, 
    0, 0, 0, 2, 1, 0, 18, 2, 2 ;

 Dg_Suspect_ice = _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, 42, _ ;

 Dg_af_fov = _, 160, 165, _, 148, _, 163, _, 169, 160, _, _, 163, 162, _, _, 
    156, 141, _, _, 153, _, _, _, 167, 48, _, 146, 162, 26, _, _, _, _, _, _, 
    _, _, 173, _, 150, 145, _, 171, _, 159, _, 162, _, 158 ;

 Dg_border_fov = 14, 46, 14, 12, 28, _, 16, _, 27, 29, 10, _, 26, 14, 2, 11, 
    17, 28, 8, 6, 25, 9, 11, 11, 44, 27, 9, 28, 16, 83, 10, 8, 9, 11, _, _, 
    _, 2, 33, 10, 32, 32, _, 50, 9, 16, 10, 32, 10, 31 ;

 Dg_chi2_Acard = 365, 710, 582, 313, 126, _, _, _, 122, 108, 113, _, 90, 109, 
    _, _, 93, 106, 84, _, 99, 99, 103, _, 97, 114, 113, 140, 114, 172, 111, 
    161, _, 74, _, _, _, _, 114, 111, 108, _, _, 89, 76, 107, 89, 98, _, _ ;

 Dg_chi2_P_Acard = 1000, 1000, 1000, 1000, 992, _, _, _, 990, 821, 786, _, 
    129, 845, _, _, 235, 752, 247, _, 462, 501, 590, _, 383, 916, 758, 999, 
    942, 999, 727, 997, _, 167, _, _, _, _, 928, 709, 792, _, _, 126, 149, 
    794, 346, 428, _, _ ;

 Dg_chi2_P_corr = _, _, _, _, 980, _, _, _, 987, 760, 750, _, 107, 765, _, _, 
    186, 714, 210, _, 428, 453, 519, _, 325, 895, 678, 999, 920, 999, 684, 
    996, _, 111, _, _, _, _, 756, 669, 687, _, _, 87, 120, 767, 302, _, _, _ ;

 Dg_chi2_P_uncorr = _, _, _, _, 985, _, _, _, 995, 730, 768, _, 170, 781, _, 
    _, 186, 742, 192, _, 437, 447, 522, _, 324, 898, 678, 999, 975, 1000, 
    653, 999, _, 160, _, _, _, _, 993, 908, 865, _, _, 80, 106, 801, 308, _, 
    _, _ ;

 Dg_chi2_corr = _, _, _, _, 121, _, _, _, 122, 106, 111, _, 89, 106, _, _, 
    92, 105, 81, _, 98, 97, 100, _, 95, 113, 108, 139, 113, 171, 108, 158, _, 
    69, _, _, _, _, 106, 109, 104, _, _, 87, 73, 106, 86, _, _, _ ;

 Dg_chi2_uncorr = _, _, _, _, 123, _, _, _, 125, 105, 112, _, 91, 107, _, _, 
    92, 106, 80, _, 98, 97, 100, _, 95, 113, 108, 139, 118, 200, 107, 180, _, 
    74, _, _, _, _, 125, 132, 110, _, _, 87, 72, 108, 87, _, _, _ ;

 Dg_galactic_Noise_Error = _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _ ;

 Dg_moonglint = _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _ ;

 Dg_num_iter_Acard = 5, 8, 8, 5, 7, _, _, _, 6, 7, 6, _, 7, 7, _, _, 7, 7, 6, 
    _, 7, 6, 7, _, 7, 7, 6, 7, 7, 7, 6, 6, _, 7, _, _, _, _, 7, 6, 7, _, _, 
    7, 6, 7, 6, 7, _, _ ;

 Dg_num_iter_corr = _, _, _, _, 20, _, _, _, 3, 20, 2, _, 2, 3, _, _, 2, 2, 
    2, _, 2, 3, 2, _, 2, 2, 3, 3, 3, 2, 2, 2, _, 2, _, _, _, _, 3, 2, 8, _, 
    _, 3, 2, 3, 2, _, _, _ ;

 Dg_num_iter_uncorr = _, _, _, _, 20, _, _, _, 3, 17, 3, _, 3, 3, _, _, 2, 2, 
    2, _, 2, 3, 3, _, 2, 2, 3, 3, 3, 3, 2, 3, _, 2, _, _, _, _, 15, 3, 8, _, 
    _, 2, 3, 3, 2, _, _, _ ;

 Dg_num_meas_l1c = 87, 220, 225, 81, 226, _, 223, _, 234, 234, 61, _, 235, 
    222, 2, 21, 216, 230, 37, 12, 235, 59, 62, 17, 225, 221, 51, 229, 222, 
    177, 48, 50, 24, 64, _, _, _, 2, 234, 38, 240, 237, _, 231, 36, 219, 36, 
    222, 63, 249 ;

 Dg_num_meas_valid = 70, 143, 190, 69, 155, _, 160, _, 182, 180, 51, _, 182, 
    191, _, 10, 182, 171, 29, 6, 181, 50, 51, 6, 163, 147, 42, 165, 189, 87, 
    38, 42, 15, 21, _, _, _, _, 171, 28, 169, 166, _, 160, 27, 183, 26, 134, 
    53, 72 ;

 Dg_quality_SSS_anom = 0, 0, 0, 0, _, 0, 0, 0, _, _, 321, 0, 151, 97, 0, 0, 
    58, 103, 369, 0, 91, 190, 178, 0, 66, 133, 177, _, 59, _, 185, _, 0, 156, 
    0, 0, 0, 0, 147, 406, 202, 0, 0, 145, 411, 186, 432, 0, 0, 0 ;

 Dg_quality_SSS_corr = _, _, _, _, _, _, _, _, _, _, 321, _, 151, 97, _, _, 
    58, 103, 369, _, 91, 190, 178, _, 66, 133, 177, _, 59, _, 185, _, _, 156, 
    _, _, _, _, 147, 406, 202, _, _, 145, 411, 186, 432, _, _, _ ;

 Dg_quality_SSS_uncorr = _, _, _, _, _, _, _, _, _, 147, 321, _, 151, 97, _, 
    _, 58, 103, 369, _, 91, 190, 178, _, 66, 133, 177, _, _, _, 185, _, _, 
    156, _, _, _, _, _, 406, 202, _, _, 145, 411, 186, 432, _, _, _ ;

 Dg_sky = 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 36, 0, 0, 0, 0, 0, 0, 0, 0, 13, 38, 34, 0, 0, 0, 0, 
    0, 0, 0, 0, 0 ;

 Dg_sun_glint_L2 = _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _ ;

 Dg_sun_glint_area = 80, 6, _, 75, _, _, _, _, 6, _, _, _, 6, _, 2, _, _, _, 
    37, _, _, 42, _, _, _, _, 27, _, _, _, 16, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _ ;

 Dg_sun_glint_fov = _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _ ;

 Dg_sun_tails = 18, 17, 31, 18, 147, _, 18, _, 15, 154, 6, _, 17, 17, _, _, 
    16, 90, 20, _, 106, 18, _, _, 103, _, 14, 16, 15, _, 7, _, _, _, _, _, _, 
    _, 172, _, 42, 58, _, 42, _, 22, _, 38, _, 84 ;

 Equiv_ftprt_diam = 46.97908, 49.76162, 48.44484, 47.27116, 51.22816, _, 
    48.11411, _, 50.61799, 51.00514, 48.98641, _, 50.90693, 47.9198, 
    64.83355, 58.7957, 48.82625, 52.60048, 54.35325, 57.81688, 51.52447, 
    49.11769, 48.67284, 59.76452, 48.73295, 58.69532, 50.39048, 54.49858, 
    47.70457, 59.14614, 51.04953, 50.18056, 57.10167, 47.11874, _, _, _, 
    65.22234, 50.3494, 54.97495, 55.26436, 55.33012, _, 49.99406, 55.67471, 
    49.46726, 56.09352, 49.15183, 50.31537, 53.96429 ;

 Grid_Point_ID = 814, 16230, 4090593, 9022, 25491, 24410, 44970, 55759, 
    74697, 81901, 63462, 88516, 1005407, 1017195, 117218, 1025437, 1038163, 
    1054563, 1019696, 1056646, 1075536, 1045794, 1078630, 1087347, 1103675, 
    1120583, 1082124, 1118994, 1130784, 1154363, 1113342, 1150794, 1159504, 
    1168188, 1156339, 1204537, 6038569, 6050362, 6078996, 6072884, 6104611, 
    6102523, 6079460, 6123532, 6094306, 6144022, 6115817, 6164506, 6159938, 
    6191161 ;

 Latitude = 84.474, 78.565, 80.915, 83.111, 73.501, 79.885, 70.735, 65.941, 
    65.152, 61.056, 62.966, 64.077, 54.48, 51.965, 58.16, 52.04, 44.882, 
    41.405, 47.555, 42.764, 34.273, 39.361, 34.868, 33.277, 25.069, 21.339, 
    27.478, 17.874, 15.737, 11.326, 17.875, 13.369, 11.428, 7.632, 5.515, 
    -2.752, -34.284, -36.546, -46.33, -43.07, -52.243, -53.147, -48.236, 
    -57.728, -51.938, -62.353, -56.375, -66.741, -65.027, -72.948 ;

 Longitude = 9.96, -8.663, 37.312, -6.626, -11.137, -24.17, -24.798, -22.766, 
    -34.694, -30.459, -22.517, -43.089, -41.245, -39.034, -48.497, -29.708, 
    -43.222, -40.729, -49.166, -35.266, -43.463, -50.001, -40.397, -38.988, 
    -47.2, -46.025, -52.93, -52.654, -51.112, -48.234, -55.05, -46.347, 
    -45.804, -48.366, -56.817, -49.091, -56.971, -54.812, -64.263, -57.778, 
    -64.657, -73.448, -74.111, -73.724, -77.577, -76.082, -81.111, -81.496, 
    -66.299, -79.85 ;

 Mean_acq_time = 7851.884, 7851.884, 7851.883, 7851.884, 7851.885, _, 
    7851.886, _, 7851.887, 7851.888, 7851.888, _, 7851.89, 7851.89, 7851.89, 
    7851.89, 7851.892, 7851.892, 7851.892, 7851.892, 7851.894, 7851.893, 
    7851.894, 7851.894, 7851.895, 7851.896, 7851.896, 7851.896, 7851.897, 
    7851.897, 7851.897, 7851.898, 7851.898, 7851.899, _, _, _, 7851.907, 
    7851.909, 7851.909, 7851.91, 7851.911, _, 7851.912, 7851.911, 7851.913, 
    7851.912, 7851.914, 7851.913, 7851.915 ;

 SSS_anom = _, _, _, _, -3.089294, _, _, _, -7.678577, -1.243866, _, _, 
    -0.4689827, -1.54398, _, _, 1.199913, 0.3051834, _, _, 0.5411835, _, _, 
    _, 0.6532974, 0.1702957, _, -0.4499054, -0.1914406, -2.226696, _, _, _, 
    _, _, _, _, _, 0.5213833, _, 1.174973, _, _, 2.259945, _, 0.3745079, _, 
    _, _, _ ;

 SSS_climatology = 65535, 65535, 65535, 65535, 2845, 65535, 65535, 65535, 
    3272, 3238, 65535, 65535, 3399, 3388, 65535, 65535, 3516, 3635, 65535, 
    65535, 3704, 65535, 65535, 65535, 3775, 3725, 65535, 3611, 3647, 3519, 
    65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 3096, 65535, 
    3089, 65535, 65535, 3519, 65535, 3317, 65535, 65535, 65535, 65535 ;

 SSS_corr = _, _, _, _, 25.62033, _, _, _, 24.53318, 33.84064, 32.24722, _, 
    33.95403, 32.52054, _, _, 36.40296, 36.42946, 33.1171, _, 37.57076, 
    35.8894, 37.47202, _, 38.40047, 37.43526, 37.26958, 35.68861, 36.15342, 
    33.87375, 33.28657, 37.18805, _, 36.11375, _, _, _, _, 34.72534, 
    36.53983, 35.23218, _, _, 36.39228, 29.04665, 34.17802, 31.0801, _, _, _ ;

 SSS_uncorr = _, _, _, _, 25.35771, _, _, _, 25.03742, 31.14113, 27.53278, _, 
    33.52202, 32.33202, _, _, 36.35791, 36.65818, 32.80346, _, 37.58318, 
    35.87761, 37.53548, _, 38.4003, 37.4213, 37.26863, 35.66409, 36.28256, 
    32.9593, 33.06751, 34.77792, _, 37.42514, _, _, _, _, 31.47838, 29.96474, 
    32.06297, _, _, 37.44894, 21.3534, 33.54051, 31.13237, _, _, _ ;

 SST = _, _, _, _, 2.188019, _, _, _, 1.405334, 9.277222, 9.560852, _, 
    8.031403, 9.728241, _, _, 17.98907, 20.44608, 8.177246, _, 25.49045, 
    22.55124, 24.41672, _, 26.38861, 26.28226, 28.05515, 26.85501, 27.04086, 
    27.36554, 27.19827, 26.45358, _, 28.6333, _, _, _, _, 8.878357, 7.94574, 
    7.01532, _, _, 5.179047, 6.895508, 1.490234, 5.518555, _, _, _ ;

 Science_Flags_Acard = 2109849, 2232729, 2109851, 2109851, 70025, 4206976, 
    12314, 4208896, 39307, 71937, 71939, 4208896, 39297, 14721, 71937, 40321, 
    16257, 16257, 69889, 73473, 39809, 40833, 40833, 39809, 68353, 11137, 
    72449, 15233, 15233, 15233, 15233, 15233, 39809, 23297, 4209152, 4203008, 
    4203520, 267523, 69891, 39041, 69889, 4329858, 4206592, 22913, 36995, 
    12417, 14721, 69913, 266666, 4329882 ;

 Science_Flags_anom = 12697, 135577, 12699, 12699, 70025, 4206976, 12314, 
    4208896, 39307, 71937, 71939, 4208896, 39297, 14721, 71937, 40321, 16257, 
    16257, 69889, 73473, 39809, 40833, 40833, 39809, 68353, 11137, 72449, 
    15233, 15233, 15233, 15233, 15233, 39809, 23297, 4209152, 4203008, 
    4203520, 267523, 69891, 39041, 69889, 4329858, 4206592, 22913, 36995, 
    12417, 14721, 69913, 266666, 4329882 ;

 Science_Flags_corr = 12697, 135577, 12699, 12699, 70025, 4206976, 12314, 
    4208896, 39307, 71937, 71939, 4208896, 39297, 14721, 71937, 40321, 16257, 
    16257, 69889, 73473, 39809, 40833, 40833, 39809, 68353, 11137, 72449, 
    15233, 15233, 15233, 15233, 15233, 39809, 23297, 4209152, 4203008, 
    4203520, 267523, 69891, 39041, 69889, 4329858, 4206592, 22913, 36995, 
    12417, 14721, 69913, 266666, 4329882 ;

 Science_Flags_uncorr = 12697, 135577, 12699, 12699, 70025, 4206976, 12314, 
    4208896, 39307, 71937, 71939, 4208896, 39297, 14721, 71937, 40321, 16257, 
    16257, 69889, 73473, 39809, 40833, 40833, 39809, 68353, 11137, 72449, 
    15233, 15233, 15233, 15233, 15233, 39809, 23297, 4209152, 4203008, 
    4203520, 267523, 69891, 39041, 69889, 4329858, 4206592, 22913, 36995, 
    12417, 14721, 69913, 266666, 4329882 ;

 Sigma_Acard = _, _, _, _, 0.6414467, _, _, _, 0.6073118, 0.5970353, 
    0.9842229, _, 0.5746502, 0.5701323, _, _, 0.5957432, 0.6526763, 1.416423, 
    _, 0.6578674, 1.159307, 1.079815, _, 0.6553078, 0.7392487, 1.40843, 
    0.8093659, 0.6887774, 1.029835, 1.40911, 1.577927, _, 1.531075, _, _, _, 
    _, 0.6233149, 1.547258, 0.6134786, _, _, 0.5567054, 1.308162, 0.5669218, 
    1.350594, _, _, _ ;

 Sigma_SSS_anom = _, _, _, _, 2.324003, _, _, _, 3.132885, 0.966469, 2.02868, 
    _, 1.135815, 0.9430208, _, _, 0.880279, 0.8424814, 3.603568, _, 
    0.7372941, 1.410482, 1.389262, _, 0.5110192, 0.8288953, 1.179508, 
    0.7761204, 0.5910576, 1.184564, 1.412123, 1.708509, _, 1.38097, _, _, _, 
    _, 0.9880466, 3.619019, 1.090589, _, _, 1.66999, 3.899885, 2.849992, 
    4.071067, _, _, _ ;

 Sigma_SSS_corr = _, _, _, _, 2.324003, _, _, _, 3.132885, 0.966469, 2.02868, 
    _, 1.135815, 0.9430208, _, _, 0.880279, 0.8424814, 3.603568, _, 
    0.7372941, 1.410482, 1.389262, _, 0.5110192, 0.8288953, 1.179508, 
    0.7761204, 0.5910576, 1.184564, 1.412123, 1.708509, _, 1.38097, _, _, _, 
    _, 0.9880466, 3.619019, 1.090589, _, _, 1.66999, 3.899885, 2.849992, 
    4.071067, _, _, _ ;

 Sigma_SSS_uncorr = _, _, _, _, 2.363697, _, _, _, 3.255715, 1.037909, 
    2.218864, _, 1.237838, 0.9506618, _, _, 0.9416327, 0.847591, 3.631229, _, 
    0.7373694, 1.410687, 1.390496, _, 0.5110149, 0.8293273, 1.179539, 
    0.7755325, 0.6068746, 1.267809, 1.397233, 1.774594, _, 1.403963, _, _, _, 
    _, 1.392263, 4.246368, 1.221886, _, _, 1.644628, 4.748276, 2.696102, 
    4.066112, _, _, _ ;

 Sigma_Tb_42_5H = _, _, _, _, 0.577449, _, _, _, 0.7016248, 0.4357364, 
    0.7184324, _, 0.5182294, 0.4466445, _, _, 0.6127065, 0.6510348, 1.078594, 
    _, 0.6280346, 0.8463717, 0.9672686, _, 0.4522795, 0.6861773, 0.771464, 
    0.6310234, 0.5428518, 0.8603384, 0.9699873, 1.077407, _, 0.8969938, _, _, 
    _, _, 0.5258167, 1.175202, 0.4580067, _, _, 0.7070469, 1.183237, 
    0.9449836, 1.146152, _, _, _ ;

 Sigma_Tb_42_5V = _, _, _, _, 0.6766798, _, _, _, 0.836141, 0.4340073, 
    0.867321, _, 0.5204526, 0.4523531, _, _, 0.6279806, 0.6525238, 1.420577, 
    _, 0.6467561, 1.009799, 1.111406, _, 0.4285015, 0.7244281, 0.9315772, 
    0.6732657, 0.5327402, 0.994175, 1.175651, 1.345838, _, 1.10738, _, _, _, 
    _, 0.4410779, 1.498369, 0.4415781, _, _, 0.7232178, 1.475247, 1.005942, 
    1.431325, _, _, _ ;

 Sigma_Tb_42_5X = _, _, _, _, 0.6028895, _, _, _, 0.7227553, 0.4707647, 
    1.148602, _, 0.5434333, 0.4466426, _, _, 0.6093559, 0.724571, 1.534314, 
    _, 0.735884, 1.209185, 1.488259, _, 0.5127047, 1.17153, 1.182312, 
    0.8735232, 0.5721648, 1.247839, 1.361563, 1.639528, _, 1.294894, _, _, _, 
    _, 0.5229029, 1.469253, 0.4604947, _, _, 0.7026207, 1.524598, 0.9363263, 
    1.502561, _, _, _ ;

 Sigma_Tb_42_5Y = _, _, _, _, 0.6898342, _, _, _, 0.8351544, 0.4710595, 
    1.162205, _, 0.5466444, 0.4519382, _, _, 0.6248335, 0.7215611, 1.384269, 
    _, 0.7465639, 1.205847, 1.498234, _, 0.4951575, 1.189994, 1.171882, 
    0.8895527, 0.5626543, 1.296721, 1.325419, 1.614335, _, 1.332812, _, _, _, 
    _, 0.4403685, 1.308366, 0.4508263, _, _, 0.7184046, 1.371611, 0.9960318, 
    1.348236, _, _, _ ;

 Sigma_WS_corr = 2785, 2591, 2602, 2800, 2577, 2813, 2811, 2657, 2590, 2476, 
    2812, 2802, 2569, 2516, 2804, 2810, 2512, 2564, 2795, 2819, 2531, 2796, 
    2806, 2803, 2501, 2571, 2809, 2563, 2492, 2773, 2814, 2811, 2805, 2813, 
    2819, 2822, 2809, 2800, 2497, 2817, 2591, 2762, 2638, 2537, 2815, 2442, 
    2817, 2233, 2788, 2810 ;

 Tb_42_5H = _, _, _, _, 78.79262, _, _, _, 79.51479, 77.55651, 78.7409, _, 
    78.34685, 78.70938, _, _, 78.59395, 78.08981, 77.98923, _, 77.24751, 
    77.54582, 77.88909, _, 75.56124, 77.1545, 75.23747, 77.5805, 77.07239, 
    78.85461, 79.09518, 77.5706, _, 76.41844, _, _, _, _, 77.31783, 82.15441, 
    77.4789, _, _, 78.97094, 81.7303, 80.2152, 80.62939, _, _, _ ;

 Tb_42_5V = _, _, _, _, 122.8353, _, _, _, 123.1669, 121.8039, 122.7644, _, 
    121.8456, 122.6062, _, _, 121.9089, 121.5505, 121.9419, _, 120.4008, 
    121.3838, 120.9691, _, 118.9925, 120.368, 119.2856, 121.3258, 120.7934, 
    122.9207, 123.3359, 120.7801, _, 120.5352, _, _, _, _, 121.3705, 
    124.1908, 121.0917, _, _, 121.4744, 125.0059, 122.3547, 123.7802, _, _, _ ;

 Tb_42_5X = _, _, _, _, 83.6256, _, _, _, 83.91153, 82.24252, 100.3814, _, 
    83.27042, 80.82545, _, _, 80.71564, 84.29158, 113.1559, _, 83.14248, 
    100.7302, 98.909, _, 78.21357, 87.19759, 100.8278, 85.83729, 79.33548, 
    91.74292, 107.2765, 103.2546, _, 95.55705, _, _, _, _, 81.20382, 
    115.7534, 85.5455, _, _, 81.94858, 117.3388, 82.30018, 116.9097, _, _, _ ;

 Tb_42_5Y = _, _, _, _, 121.2638, _, _, _, 122.1012, 120.5553, 104.5532, _, 
    120.3218, 123.8646, _, _, 123.1848, 118.7413, 90.19884, _, 117.9917, 
    101.6551, 103.4226, _, 119.8658, 113.808, 97.22634, 116.5288, 121.9944, 
    113.4571, 98.57793, 98.55373, _, 104.8676, _, _, _, _, 120.8139, 
    93.92569, 116.349, _, _, 121.7193, 92.58741, 123.3886, 90.66586, _, _, _ ;

 WS = _, _, _, _, 9.118509, _, _, _, 8.506406, 5.581868, 5.255404, _, 
    7.568759, 7.81521, _, _, 9.663113, 10.00159, 4.873579, _, 10.20495, 
    8.297751, 10.58992, _, 6.278353, 8.653219, 3.985853, 10.02652, 9.747353, 
    9.001951, 10.41351, 10.25866, _, 3.515022, _, _, _, _, 3.135072, 
    12.05383, 3.885997, _, _, 9.806511, 12.50787, 14.0133, 11.63738, _, _, _ ;

 WS_corr = 11325, 9247, 4399, 10719, 4535, 12061, 8988, 9968, 7914, 2663, 
    5241, 4169, 7537, 6487, 6868, 6138, 10902, 9537, 4748, 4534, 9829, 7710, 
    11034, 7867, 5300, 9102, 3165, 8717, 7441, 8478, 9979, 9683, 8045, 3670, 
    3140, 4622, 11455, 12895, 2708, 12218, 4120, 15710, 5772, 11975, 12639, 
    15145, 11676, 1850, 16455, 9713 ;

 X_swath = -414.0223, -113.8237, 72.9677, -424.9457, 199.7495, _, _, _, 
    -169.8757, 190.8608, 471.225, _, -185.8288, 31.19449, _, 629.5717, 
    -60.22084, 236.2844, -569.8598, _, 214.5479, -477.9211, 467.9586, 
    643.6125, 110.6364, 324.5805, -504.4055, -268.7122, -58.32698, 353.2138, 
    -517.254, 501.2082, 609.0753, 431.5117, _, _, _, _, 143.988, 575.2241, 
    267.69, _, _, -117.7976, -583.241, -60.96313, -588.8839, -105.4338, _, _ ;
}
