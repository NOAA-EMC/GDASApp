netcdf sst.nc {
dimensions:
	Location = 201 ;
	nvars = 1 ;
variables:
	int Location(Location) ;
		Location:suggested_chunk_dim = 201LL ;
	float nvars(nvars) ;
		nvars:suggested_chunk_dim = 100LL ;

// global attributes:
		string :_ioda_layout = "ObsGroup" ;
		:_ioda_layout_version = 0 ;
		:nrecs = 1 ;
		:converter = "gds2_sst2ioda.py" ;
		:processing_level = "L3U" ;
		:nvars = 1 ;
		:date_time = 2018041512 ;
		:nlocs = 201 ;
		:nobs = 201 ;
		:thinning = 0.99999 ;
		:sensor = "AVHRR_GAC" ;
		:platform = "NOAA-19" ;
data:

 Location = 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 nvars = 0 ;

group: MetaData {
  variables:
  	int64 dateTime(Location) ;
  		dateTime:_FillValue = -3732782400LL ;
  		string dateTime:units = "seconds since 2018-04-15T12:00:00Z" ;
  	string date_time(Location) ;
  		string date_time:_FillValue = "" ;
  	float latitude(Location) ;
  		latitude:_FillValue = 9.96921e+36f ;
  	float longitude(Location) ;
  		longitude:_FillValue = 9.96921e+36f ;
  	string variable_names(nvars) ;
  		string variable_names:_FillValue = "" ;
  data:

   dateTime = -40813, -41195, -41918, -41960, -42007, -42014, -42017, -36233,
      -34897, -33232, -35478, -35689, -35678, -35735, -35715, -35743, -35785,
      -35793, -35785, -35883, -35908, -29089, -29166, -29200, -29259, -29550,
      -29582, -29905, -30064, -32128, -31982, -26780, -26555, -26398, -26400,
      -26190, -26095, -25842, -25787, -22996, -23045, -23068, -23191, -23338,
      -23439, -23523, -23903, -23962, -21107, -21068, -20959, -20775, -20786,
      -20717, -20347, -19585, -14862, -14722, -16968, -17083, -17174, -17163,
      -17576, -17598, -17587, -10919, -11331, -11437, -11469, -8438, -8172,
      -8145, -7703, -7664, -7472, -7230, -3743, -3867, -4812, -5357, -5363,
      -2328, -2212, -2116, -1825, -1820, -1681, -1671, -1683, -1682, -1564,
      2231, 3179, 870, 826, 3842, 3926, 3954, 4056, 4074, 4194, 4243, 4264,
      4388, 4518, 9214, 9281, 10234, 10274, 10252, 10296, 10590, 10635,
      10608, 10667, 14008, 13880, 13869, 13773, 13199, 12874, 12817, 12636,
      12659, 10827, 12394, 15350, 15513, 15596, 16616, 16664, 16851, 17139,
      17170, 20450, 20414, 20423, 19972, 19922, 19871, 19825, 19825, 19635,
      19398, 19281, 19262, 19225, 19178, 19013, 18943, 18893, 18909, 18263,
      21885, 22125, 22658, 22794, 24800, 27876, 25968, 25956, 28112, 28166,
      25762, 28718, 32111, 32144, 32008, 31987, 31902, 31528, 28826, 28868,
      30927, 30882, 34355, 34414, 34928, 34986, 35036, 35499, 38222, 38147,
      38096, 37996, 37982, 37870, 37785, 37711, 37597, 37596, 37539, 37510,
      36943, 40469, 40520, 40518, 41066, 41181, 41548, 41722 ;

   latitude = 58.91, 36.77, -5.189998, -8.749998, -9.209998, -11.37, -12.21,
      -30.81, 44.97, 31.83, 12.69, 1.890002, 1.550002, -0.449998, -1.009998,
      -1.069998, -3.889998, -4.049998, -5.009998, -9.989998, -11.23, 27.99,
      25.07, 21.37, 18.37, 0.430002, -0.689998, -19.11, -28.89, -30.09,
      -37.57, 15.45, -0.02999799, -7.609998, -8.089998, -21.83, -25.87,
      -41.25, -44.51, 28.63, 24.47, 21.53, 17.03, 5.910002, 0.330002,
      -3.189998, -24.83, -27.81, 40.85, 37.27, 32.95, 21.43, 20.71, 17.75,
      -5.669998, -47.19, 31.81, 23.51, 23.27, 16.43, 9.950002, 9.130002,
      -12.39, -13.63, -15.51, 16.33, -4.809998, -10.91, -13.17, 14.95,
      -0.669998, -1.689998, -28.69, -30.87, -40.93, -56.17, 75.23, 69.91,
      15.65, -14.41, -15.29, 16.13, 10.39, 2.850002, -13.75, -14.19, -20.07,
      -21.29, -22.25, -22.33, -28.95, 66.39, 53.09, -9.149998, -11.75, 13.47,
      8.850002, 6.530002, 0.930002, -0.149998, -7.929998, -10.55, -11.01,
      -19.73, -27.47, 56.17, 51.93, -2.429998, -4.749998, -5.109998,
      -5.869998, -23.33, -24.47, -24.79, -26.97, 42.07, 36.67, 36.01, 28.47,
      -3.769998, -21.71, -25.51, -35.57, -35.81, -37.35, -50.17, 55.21,
      47.49, 41.33, -17.57, -21.37, -31.09, -47.69, -50.07, 62.31, 60.27,
      59.67, 35.89, 32.99, 30.05, 26.29, 25.37, 16.09, 1.590002, -5.749998,
      -6.289998, -10.31, -12.45, -20.11, -24.85, -26.97, -26.99, -63.71,
      31.59, 17.41, -13.87, -22.57, -41.61, 39.39, 27.23, 24.99, 23.49,
      21.55, 13.71, -10.79, 29.19, 28.51, 23.43, 22.27, 17.45, -7.489998,
      -16.65, -17.43, -39.65, -42.59, 19.69, 15.79, -14.25, -17.41, -22.57,
      -47.19, 27.01, 25.01, 20.03, 15.27, 13.89, 6.230002, 3.550002,
      -1.489998, -8.429997, -8.469997, -10.93, -12.59, -45.69, 19.47, 16.73,
      16.69, -16.89, -20.33, -42.73, -54.77 ;

   longitude = -146.77, -138.63, -127.65, -134.05, -119.81, -129.79, -134.81,
      -148.69, -176.33, 31.52999, -161.01, -149.97, -155.71, -147.33,
      -157.67, -148.01, -149.67, -147.95, -156.25, -150.59, -148.97, 168.45,
      177.67, 169.21, 172.01, 170.07, 174.41, -179.27, 177.51, 1.809996,
      -5.130004, -17.29, -3.950004, -16.79, -12.55, -3.790004, -17.27,
      -15.91, -15.99, 156.91, 148.61, 141.31, 157.43, 144.53, 147.39, 156.53,
      164.27, 167.61, -30.03, -22.47, -40.95, -34.53, -26.09, -33.51, -26.81,
      -56.07, -46.83, -47.95, 132.81, 133.65, 126.99, 118.89, 138.61, 139.15,
      122.17, 92.50999, 113.47, 115.09, 113.71, -80.95, -83.95, -88.07,
      -84.49001, -85.51, -98.15, -84.15, 25.67, 42.94999, 67.81, 84.34999,
      81.09, -109.67, -118.61, -106.95, -113.31, -112.51, -127.25, -124.17,
      -113.89, -113.63, -116.77, 10.91, -140.25, 52.02999, 52.39, -136.85,
      -139.79, -136.03, -139.51, -139.85, -136.21, -138.79, -143.83, -135.37,
      -134.95, -143.37, -143.01, -165.79, -166.51, -155.11, -168.03, -170.13,
      -178.57, -167.83, -176.11, -15.97, -3.190004, -3.130004, -11.81,
      1.829996, 11.89, 10.11, 15.29, 3.549996, -172.33, 15.91, -168.73,
      174.71, -176.05, 164.31, 170.67, 159.81, 154.63, 157.43, -40.59,
      -39.29, -46.19, -19.45, -18.89, -18.31, -26.91, -31.93, -18.51, -19.89,
      -21.11, -17.79, -29.09, -24.25, -10.85, -13.43, -8.810004, -13.93,
      2.669996, 155.27, 152.85, 145.99, 151.13, -45.35, 130.49, -54.45,
      -62.13, 137.37, 131.07, -59.69, 125.01, -75.91, -90.23, -72.83,
      -72.35001, -70.21, -85.07, 120.31, 109.17, -59.59, -60.53, 90.78999,
      93.46999, 86.74999, 84.73, 100.71, 76.38999, -110.47, -93.75, -107.01,
      -99.67, -102.53, -107.39, -93.09, -96.47, -96.41, -96.37, -90.85,
      -90.49001, -82.77, 70.41, 67.73, 69.17, 72.31, 51.64999, 50.84999, 61.07 ;

   variable_names = "sea_surface_temperature" ;
  } // group MetaData

group: ObsError {
  variables:
  	float seaSurfaceTemperature(Location) ;
  		seaSurfaceTemperature:_FillValue = 9.96921e+36f ;
  data:

   seaSurfaceTemperature = 0.29, 0.29, 0.39, 0.47, 0.39, 0.39, 0.42, 0.37,
      0.32, 0.39, 0.39, 0.4, 0.39, 0.42, 0.39, 0.39, 0.34, 0.37, 0.39, 0.48,
      0.48, 0.29, 0.27, 0.33, 0.43, 0.48, 0.58, 0.39, 0.36, 0.22, 0.28, 0.4,
      0.54, 0.28, 0.29, 0.32, 0.24, 0.27, 0.28, 0.29, 0.32, 0.42, 0.43, 0.48,
      0.63, 0.48, 0.32, 0.36, 0.27, 0.26, 0.31, 0.36, 0.26, 0.21, 0.25, 0.29,
      0.23, 0.24, 0.37, 0.39, 0.44, 0.52, 0.48, 0.48, 0.48, 0.53, 0.56, 0.51,
      0.45, 0.34, 0.3, 0.19, 0.24, 0.29, 0.27, 0.42, 0.33, 0.33, 0.53, 0.39,
      0.41, 0.23, 0.33, 0.29, 0.19, 0.25, 0.34, 0.36, 0.19, 0.21, 0.27, 0.39,
      0.29, 0.44, 0.48, 0.32, 0.48, 0.39, 0.27, 0.17, 0.2, 0.41, 0.26, 0.44,
      0.32, 0.28, 0.28, 0.29, 0.3, 0.33, 0.46, 0.14, 0.34, 0.22, 0.34, 0.29,
      0.29, 0.29, 0.43, 0.48, 0.29, 0.29, 0.28, 0.31, 0.25, 0.28, 0.28, 0.33,
      0.29, 0.42, 0.27, 0.31, 0.27, 0.28, 0.32, 0.28, 0.29, 0.36, 0.34, 0.45,
      0.29, 0.35, 0.34, 0.48, 0.45, 0.45, 0.46, 0.39, 0.33, 0.32, 0.35, 0.3,
      0.3, 0.24, 0.3, 0.22, 0.27, 0.3, 0.28, 0.3, 0.39, 0.27, 0.33, 0.52,
      0.22, 0.29, 0.36, 0.36, 0.42, 0.48, 0.48, 0.46, 0.53, 0.27, 0.29, 0.52,
      0.49, 0.26, 0.23, 0.34, 0.32, 0.44, 0.38, 0.44, 0.48, 0.48, 0.52, 0.5,
      0.35, 0.31, 0.31, 0.39, 0.36, 0.29, 0.51, 0.45, 0.5, 0.3, 0.32, 0.27,
      0.21 ;
  } // group ObsError

group: ObsValue {
  variables:
  	float seaSurfaceTemperature(Location) ;
  		seaSurfaceTemperature:_FillValue = 9.96921e+36f ;
  data:

   seaSurfaceTemperature = 5.803994, 13.77201, 27.064, 27.87, 26.804, 27.56,
      28.04401, 23.72399, 5.648, 18.796, 27.22001, 27.57401, 27.27401,
      26.31599, 26.88601, 26.71201, 27.69399, 27.76599, 27.99201, 29.282,
      29.158, 20.49, 22.51001, 25.30799, 26.21601, 29.93198, 28.80801,
      27.218, 23.48199, 21.332, 17.88, 18.09201, 28.69399, 28.20799,
      27.52001, 23.73, 25.448, 16.22801, 11.512, 19.95001, 25.152, 25.94599,
      27.108, 30.13799, 30.17001, 30.59599, 25.03801, 23.708, 15.966,
      17.34999, 20.70201, 22.19199, 20.86601, 22.85399, 28.68199, 12.99401,
      21.56801, 23.868, 26.36601, 28.03, 29.3, 29.282, 30.19199, 30.42599,
      30.96801, 29.74399, 29.97799, 30.94201, 30.21599, 27.03999, 21.54199,
      24.39801, 21.08001, 21.15201, 14.18999, 6.417985, 0.9120085, 1.09599,
      29.56199, 27.56801, 27.42999, 27.35798, 27.83399, 28.49199, 25.51601,
      25.26, 26.60399, 26.15399, 25.008, 25.056, 25.03201, 6.167985,
      6.300011, 29.50001, 28.94001, 25.94, 27.66201, 27.76801, 25.988,
      26.44201, 27.26599, 28.226, 28.69601, 27.536, 25.972, 5.996015,
      5.86601, 27.63, 28.854, 27.80999, 29.11199, 26.074, 24.92398, 24.782,
      24.25601, 13.10801, 15.238, 15.362, 17.10798, 31.26999, 20.30999,
      20.714, 19.51001, 19.93201, 19.314, 4.237989, 4.211993, 3.711993,
      9.389996, 27.23799, 25.79201, 23.59601, 11.88599, 10.11001, 3.012011,
      4.411992, -1.927994, 17.23599, 18.82001, 19.76399, 21.04601, 21.82199,
      21.10999, 29.21801, 28.53401, 28.57801, 28.14401, 27.05801, 24.99401,
      25.41801, 24.67, 25.43999, 0.08600003, 19.12601, 27.44599, 28.01801,
      25.87999, 16.278, 8.505994, 24.53199, 25.18201, 24.6, 26.978, 27.11801,
      30.42799, 23.09, 22.23598, 25.93399, 26.22599, 27.09799, 25.372,
      30.39801, 27.93799, 17.91599, 15.72001, 28.846, 29.122, 27.20201,
      26.73599, 23.46399, 7.969999, 20.43399, 24.03599, 24.56201, 30.00001,
      29.84599, 29.97601, 28.97599, 26.50001, 27.156, 27.18799, 25.97801,
      25.40001, 11.42001, 28.83, 29.22801, 29.294, 27.58001, 27.64801,
      10.55799, 3.594002 ;
  } // group ObsValue

group: PreQc {
  variables:
  	float seaSurfaceTemperature(Location) ;
  		seaSurfaceTemperature:_FillValue = 9.96921e+36f ;
  data:

   seaSurfaceTemperature = 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
      0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
      0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
      0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
      0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
      0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
      0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
      0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
      0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;
  } // group PreQc
}
