netcdf sss.nc {
dimensions:
	Location = 100 ;
	nvars = 1 ;
variables:
	int Location(Location) ;
		Location:suggested_chunk_dim = 100LL ;
	float nvars(nvars) ;
		nvars:suggested_chunk_dim = 100LL ;

// global attributes:
		string :_ioda_layout = "ObsGroup" ;
		:_ioda_layout_version = 0 ;
		:nrecs = 1 ;
		:nvars = 1 ;
		:odb_version = 1LL ;
		:date_time = 2018041512 ;
		:nlocs = 100LL ;
		:nobs = 100LL ;
		:history = "Fri Apr 19 08:41:14 2019: ncks -d nlocs,1,1000000,10000 sss.orig.nc -O sst.nc" ;
		:NCO = "4.7.2" ;
data:

 Location = 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
    0, 0, 0, 0, 0, 0 ;

 nvars = 0 ;

group: MetaData {
  variables:
  	int64 dateTime(Location) ;
  		dateTime:_FillValue = -3732782400LL ;
  		string dateTime:units = "seconds since 2018-04-15T12:00:00Z" ;
  	string date_time(Location) ;
  		string date_time:_FillValue = "" ;
  	float latitude(Location) ;
  		latitude:_FillValue = 9.96921e+36f ;
  	float longitude(Location) ;
  		longitude:_FillValue = 9.96921e+36f ;
  	int sequenceNumber(Location) ;
  		sequenceNumber:_FillValue = -2147483647 ;
  	string variable_names(nvars) ;
  		string variable_names:_FillValue = "" ;
  data:

   dateTime = 16413, -15923, -37695, 14766, -25781, -11737, -9986, 20459,
      -25203, -18263, 36958, 21046, -11400, -23577, -32343, -4229, -19814,
      -19361, 9764, 22504, -19662, 1093, -37076, 22639, -38226, 38470, 3355,
      -21918, -28049, 32159, -1882, 6817, 28001, 5033, -18020, -33747, 25053,
      42188, -15155, 36241, 761, -31254, -15877, 7592, 20573, -8920, 29349,
      29808, 21036, 31289, -10162, 11895, -22210, 12609, 27289, 2940, 32325,
      -23540, 7420, 21173, -37473, 25112, -11645, -3995, 23491, -30758,
      24175, -34669, 27365, 21227, 43137, -5626, -15018, -25329, -12130,
      -12186, -32019, -16964, 12260, -19083, 2815, -31577, -11805, 27481,
      -17853, -38072, 29789, -8915, 43012, -26812, -27762, -33971, -20603,
      3250, -20704, 42063, 42910, 9413, -37307, -31455 ;

   latitude = 53.879, -58.38232, 0.393135, -46.62201, 0.3569438, 37.38496,
      -58.87528, -64.11797, 32.36138, 75.8694, -49.12336, -27.39389, 25.3784,
      39.12261, -34.36073, -50.38835, 0.884598, 28.35575, 6.134513, 63.87992,
      10.13324, -19.62038, 35.38895, 66.38779, -39.14023, -47.11112,
      -18.87907, -61.36031, -41.6361, -61.61643, 13.61734, -10.87163,
      34.38682, 72.36931, 60.62663, -60.38211, -42.64268, -6.871958,
      -64.62761, -6.131754, -2.378339, 24.61968, -61.36315, -59.37663,
      -57.13705, -50.12148, 53.11937, 34.37182, -20.87342, -59.36716,
      -57.62246, 37.1406, -34.88064, 2.888079, -8.607044, -52.12254,
      -57.8832, 37.8768, -43.11407, -12.37021, 12.12483, -38.37106, 40.37134,
      -65.13678, 58.61689, 53.35913, 9.118921, -4.877728, 3.642554,
      -18.13534, -56.38377, 27.12191, -57.11341, 32.64145, 60.38355,
      70.39142, -14.36325, 5.119036, 15.39068, 45.37792, -56.89023, 11.36977,
      41.8684, 8.370608, 50.36518, -29.38099, 28.11311, -45.87344, -49.12109,
      -63.39182, -65.10889, -44.85678, -46.86501, -30.36576, -43.63494,
      -0.8765696, -51.63343, -9.134258, 20.61064, 20.11235 ;

   longitude = 4.115798, 327.8615, 248.3797, 44.38053, 201.8728, 324.8867,
      294.0996, 17.3724, 188.1367, 43.91171, 110.8501, 10.37052, 318.6276,
      18.88903, 227.636, 279.3855, 172.6065, 165.1211, 52.86695, 330.1345,
      170.1191, 258.1304, 234.6186, 333.8995, 251.132, 297.3483, 76.89408,
      348.4011, 25.36266, 332.1636, 94.8727, 236.8727, 327.3827, 32.67982,
      355.6476, 36.36999, 154.8804, 97.62099, 179.1315, 119.6152, 270.8696,
      213.1319, 327.116, 230.1518, 18.37139, 144.6165, 160.592, 153.3711,
      8.64412, 117.3863, 304.6573, 227.6308, 354.8997, 216.3867, 338.3861,
      86.59863, 336.36, 19.87214, 237.3763, 3.612482, 241.6204, 158.8994,
      327.3783, 257.3757, 188.6524, 206.8672, 170.8689, 53.62115, 333.1209,
      4.131203, 78.86398, 294.1184, 163.8975, 187.8797, 338.088, 353.3509,
      229.1338, 340.6393, 220.6252, 157.6046, 82.86684, 217.1175, 331.1054,
      330.3774, 352.1118, 257.6353, 147.6305, 133.653, 77.65506, 223.3561,
      11.3523, 38.86535, 183.6522, 76.38167, 186.3695, 96.36871, 85.86997,
      51.61628, 238.3724, 217.1181 ;

   sequenceNumber = 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
      1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
      1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
      1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
      1, 1, 1, 1, 1, 1, 1, 1, 1 ;

   variable_names = "sea_surface_salinity" ;
  } // group MetaData

group: ObsError {
  variables:
  	float seaSurfaceSalinity(Location) ;
  		seaSurfaceSalinity:_FillValue = 9.96921e+36f ;
  data:

   seaSurfaceSalinity = 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
      1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
      1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
      1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
      1, 1, 1, 1, 1, 1, 1, 1, 1, 1 ;
  } // group ObsError

group: ObsValue {
  variables:
  	float seaSurfaceSalinity(Location) ;
  		seaSurfaceSalinity:_FillValue = 9.96921e+36f ;
  data:

   seaSurfaceSalinity = 33.71178, 34.27895, 34.89477, 33.47415, 35.26365,
      35.16874, 34.30404, 34.09843, 34.96246, 0.007955075, 35.2322, 35.57863,
      37.57914, 38.05683, 34.03303, 33.31181, 33.65787, 35.14495, 36.04657,
      34.5812, 34.02576, 36.25037, 32.16301, 34.79661, 34.63808, 33.19758,
      34.36973, 36.37263, 35.16792, 33.12465, 32.51355, 35.36753, 36.12861,
      34.40482, 35.7425, 35.411, 35.9472, 34.48295, 32.57633, 25.14996,
      34.82872, 34.71701, 35.64753, 34.48979, 34.17043, 32.8913, 0.0047155,
      35.08466, 35.65135, 32.68414, 34.3378, 33.15457, 35.72908, 34.25256,
      36.46022, 32.59492, 33.59892, 34.7174, 33.43561, 36.39915, 34.19456,
      35.34409, 36.00577, 32.72109, 31.62992, 33.06574, 33.46413, 35.41788,
      35.51361, 36.36302, 33.78024, 37.16262, 32.05506, 34.65675, 35.83234,
      34.34883, 36.18774, 33.99451, 33.84148, 32.32932, 36.14341, 33.85884,
      35.04386, 36.04567, 36.23658, 36.13433, 34.53632, 31.36066, 33.58314,
      33.99441, 35.13243, 33.27727, 35.24531, 36.08514, 35.2952, 31.50171,
      34.44715, 35.18509, 34.1835, 35.66429 ;
  } // group ObsValue

group: PreQC {
  variables:
  	int seaSurfaceSalinity(Location) ;
  		seaSurfaceSalinity:_FillValue = -2147483647 ;
  data:

   seaSurfaceSalinity = 8224, 2048, 0, 4096, 0, 0, 128, 2048, 0, 28192, 0,
      8192, 0, 8192, 0, 8192, 8192, 0, 8192, 8224, 8192, 0, 8224, 27136, 0,
      8192, 0, 2048, 0, 2048, 40960, 0, 0, 27136, 8192, 2048, 0, 0, 18432,
      9472, 0, 0, 2048, 2048, 6144, 0, 28416, 0, 8192, 2048, 2048, 0, 0, 0,
      0, 0, 2048, 8448, 0, 0, 32, 0, 32768, 18432, 14336, 0, 8192, 0, 32768,
      0, 2048, 0, 0, 0, 0, 59392, 0, 32768, 128, 2048, 2048, 32, 0, 32, 8192,
      0, 0, 4096, 128, 2048, 6144, 0, 0, 0, 0, 40960, 0, 0, 32, 0 ;
  } // group PreQC
}
