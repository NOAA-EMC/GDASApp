netcdf output_1 {
dimensions:
	Rows = 15 ;
	Columns = 45 ;
variables:
	float IceConc(Rows, Columns) ;
		IceConc:_FillValue = -999.f ;
		IceConc:coordinates = "Longitude Latitude" ;
		IceConc:long_name = "Ice Concentration" ;
		IceConc:units = "%" ;
		IceConc:valid_range = 0.f, 100.f ;
	byte IceMap(Rows, Columns) ;
		IceMap:_FillValue = -3b ;
		IceMap:coordinates = "Longitude Latitude" ;
		IceMap:long_name = "Ice Cover map codes" ;
		IceMap:units = "1" ;
		IceMap:valid_range = -2b, 2b ;
	float IceRetrPct ;
		IceRetrPct:long_name = "% of valid ice cover and concentration retrievals of all water pixels" ;
		IceRetrPct:units = "%" ;
		IceRetrPct:_FillValue = 0.f ;
		IceRetrPct:valid_range = 0.f, 100.f ;
	float IceSrfTemp(Rows, Columns) ;
		IceSrfTemp:_FillValue = -999.f ;
		IceSrfTemp:coordinates = "Longitude Latitude" ;
		IceSrfTemp:long_name = "Ice Surface Temp" ;
		IceSrfTemp:units = "Kelvin(K)" ;
		IceSrfTemp:valid_range = 100.f, 390.f ;
	float IceTermntPct ;
		IceTermntPct:long_name = "% of terminated ice cover and concentration retrievals of all processed pixels" ;
		IceTermntPct:units = "%" ;
		IceTermntPct:_FillValue = 0.f ;
		IceTermntPct:valid_range = 0.f, 100.f ;
	float Latitude(Rows, Columns) ;
		Latitude:long_name = "Latitude" ;
		Latitude:_FillValue = -999.f ;
		Latitude:units = "degrees_north" ;
		Latitude:valid_range = -90.f, 90.f ;
		Latitude:comments = "Pixel latitude in field Latitude (degree)" ;
	float Longitude(Rows, Columns) ;
		Longitude:long_name = "Longitude" ;
		Longitude:_FillValue = -999.f ;
		Longitude:units = "degrees_east" ;
		Longitude:valid_range = -180.f, 180.f ;
		Longitude:comments = "Pixel longitude in field Longitude (degree)" ;
	float MaxIceConc ;
		MaxIceConc:long_name = "Max ice concentration retrieval" ;
		MaxIceConc:_FillValue = -999.f ;
		MaxIceConc:units = "%" ;
	float MeanIceConc ;
		MeanIceConc:long_name = "Mean ice concentration retrieval" ;
		MeanIceConc:_FillValue = -999.f ;
		MeanIceConc:units = "%" ;
	float MinIceConc ;
		MinIceConc:long_name = "Min ice concentration retrieval" ;
		MinIceConc:_FillValue = -999.f ;
		MinIceConc:units = "%" ;
	byte NumOfQACategories ;
		NumOfQACategories:long_name = "Number of QA flag values" ;
		NumOfQACategories:_FillValue = -128b ;
		NumOfQACategories:units = "1" ;
	int QCFlags(Rows, Columns) ;
		QCFlags:_FillValue = -1 ;
		QCFlags:coordinates = "Longitude Latitude" ;
		QCFlags:long_name = "QCFlags" ;
		QCFlags:units = "1" ;
	float STDIceConc ;
		STDIceConc:long_name = "Standard deviation of ice concentration retrievals" ;
		STDIceConc:_FillValue = -999.f ;
		STDIceConc:units = "%" ;
	byte SearchWindowSize ;
		SearchWindowSize:long_name = "Pixel size of search window to determine tie-point" ;
		SearchWindowSize:_FillValue = -128b ;
		SearchWindowSize:units = "1" ;
	int StartColumn ;
		StartColumn:long_name = "Start column index" ;
		StartColumn:units = "1" ;
	int StartRow ;
		StartRow:long_name = "Start row index" ;
		StartRow:units = "1" ;
	byte SummaryQC_Ice_Concentration(Rows, Columns) ;
		SummaryQC_Ice_Concentration:_FillValue = -128b ;
		SummaryQC_Ice_Concentration:coordinates = "Longitude Latitude" ;
		SummaryQC_Ice_Concentration:long_name = "User-level summary QC: 0=Normal, 1=Uncertain, 2=Non-Retrievable, 3=Bad" ;
		SummaryQC_Ice_Concentration:units = "1" ;
		SummaryQC_Ice_Concentration:valid_range = 0b, 3b ;
	int TotDaytimePixs ;
		TotDaytimePixs:long_name = "Total number of daytime valid retrievals" ;
		TotDaytimePixs:_FillValue = 0 ;
		TotDaytimePixs:units = "1" ;
	int TotIceRetrvls ;
		TotIceRetrvls:long_name = "Total number of valid ice cover and concentration retrievals" ;
		TotIceRetrvls:_FillValue = 0 ;
		TotIceRetrvls:units = "1" ;
	int TotIceTermnt ;
		TotIceTermnt:long_name = "Total number of terminated ice cover and concentration retrievals" ;
		TotIceTermnt:_FillValue = 0 ;
		TotIceTermnt:units = "1" ;
	int TotNighttimePixs ;
		TotNighttimePixs:long_name = "Total number of nighttime valid retrievals" ;
		TotNighttimePixs:_FillValue = 0 ;
		TotNighttimePixs:units = "1" ;
	int TotWaterPixs ;
		TotWaterPixs:long_name = "Total number of pixels w. water surface" ;
		TotWaterPixs:_FillValue = 0 ;
		TotWaterPixs:units = "1" ;
	int Tot_QA_BadData ;
		Tot_QA_BadData:long_name = "Total number of pixels with QA category 4 (Bad data)" ;
		Tot_QA_BadData:_FillValue = 0 ;
		Tot_QA_BadData:units = "1" ;
	int Tot_QA_Nonretrievable ;
		Tot_QA_Nonretrievable:long_name = "Total number of pixels with QA category 3 (Non-retrievable)" ;
		Tot_QA_Nonretrievable:_FillValue = 0 ;
		Tot_QA_Nonretrievable:units = "1" ;
	int Tot_QA_Normal ;
		Tot_QA_Normal:long_name = "Total number of pixels with QA category 1 (Normal of optimal)" ;
		Tot_QA_Normal:_FillValue = 0 ;
		Tot_QA_Normal:units = "1" ;
	int Tot_QA_Uncertain ;
		Tot_QA_Uncertain:long_name = "Total number of pixels with QA category 2 (Uncertain or suboptimal)" ;
		Tot_QA_Uncertain:_FillValue = 0 ;
		Tot_QA_Uncertain:units = "1" ;
	int64 cloud_mask_granule_level_quality_flag ;
		cloud_mask_granule_level_quality_flag:long_name = "Cloud Mask Granule Level Degradation Quality Flag" ;
		cloud_mask_granule_level_quality_flag:flag_values = 0LL, 1LL, 63LL ;
		cloud_mask_granule_level_quality_flag:flag_meanings = "Missing_Channel_Degradation Missing_Ancillary_SST_Degradation Complete_IR_Failure" ;
		cloud_mask_granule_level_quality_flag:units = "1" ;
		cloud_mask_granule_level_quality_flag:_FillValue = -999LL ;
		cloud_mask_granule_level_quality_flag:valid_range = 0LL, 63LL ;
	ubyte quality_information ;
		quality_information:long_name = "total number of retrievals, percentage of optimal retrievals, percentage_sub_optimal_retrievals, percentage of bad retrievals" ;
		quality_information:total_number_retrievals = 2450029 ;
		quality_information:percentage_optimal_retrievals = 1.511003f ;
		quality_information:percentage_sub_optimal_retrievals = 2.04471f ;
		quality_information:percentage_bad_retrievals = 96.44428f ;

// global attributes:
		:Conventions = "CF-1.6,ACDD 1.3" ;
		:Metadata_Conventions = "CF-1.6, Unidata Dataset Discovery v1.0" ;
		:standard_name_vocabulary = "CF Standard Name Table v76" ;
		:institution = "DOC/NOAA/NESDIS/OSPO > Office of Satellite and Product Operations, NESDIS, NOAA, U.S. Department of Commerce." ;
		:naming_authority = "gov.noaa.nesdis.ncei." ;
		:processing_level = "NOAA Level 2" ;
		:production_site = "NCCF" ;
		:production_environment = "prod" ;
		:sensor_band_identifier = "M3,M5,M7,M10,M15,M16" ;
		:sensor_band_central_radiation_wavelength = "0.488um,0.672um,0.865um,1.61um,10.763um,12.013um" ;
		:satellite_name = "NOAA-20" ;
		:instrument = "VIIRS" ;
		:project = "NESDIS Common Cloud Framework" ;
		:summary = "Enterprise Ice Concentration/ Ice Mask/ Ice Surface Temperature Products" ;
		:history = "Tue Aug 20 14:14:39 2024: ncks -d Columns,1,90,2 -d Rows,1,30,2 JRR-IceConcentration_v3r3_j01_s202406181055311_e202406181056538_c202406181202563.nc output_1.ncn\nEnterprise Ice Concentration Algorithm v1.1.0" ;
		:references = "N/A" ;
		:resolution = "750M" ;
		:time_coverage_start = "2024-06-18T10:55:31Z" ;
		:time_coverage_end = "2024-06-18T10:56:53Z" ;
		:date_created = "2024-06-18T12:02:56Z" ;
		:geospatial_lat_units = "degrees_north" ;
		:geospatial_lon_units = "degrees_east" ;
		:publisher_name = "DOC/NOAA/NESDIS/OSPO > Office of Satellite and Product Operations, NESDIS, NOAA, U.S. Department of Commerce." ;
		:publisher_email = "espcoperations@noaa.gov" ;
		:publisher_url = "http://www.ospo.noaa.gov" ;
		:creator_email = "jkey@ssec.wisc.edu" ;
		:creator_name = "DOC/NOAA/NESDIS/STAR > Cryosphere Team, Center for Satellite Applications and Research, NESDIS, NOAA, U.S. Department of Commerce" ;
		:creator_url = "http://www.star.nesdis.noaa.gov" ;
		:source = "L1b data, JRR-CloudMask, JRR-CloudHeight" ;
		:keywords = "EARTH SCIENCE, CRYOSPHERE, SEA ICE, SEA ICE CONCENTRATION, ICE FRACTION, ICE EXTENT, ICE EDGES" ;
		:cdm_data_type = "Swath" ;
		:platform = "NOAA-20" ;
		:title = "JRR_IceConcentration" ;
		:metadata_link = "JRR-IceConcentration_v3r3_j01_s202406181055311_e202406181056538_c202406181202563.nc" ;
		:history_package = "Delivery Package v3r3" ;
		:product_version = "v3r3" ;
		:keywords_vocabulary = "NASA Global Change Master Directory (GCMD) Science Keywords" ;
		:geospatial_lat_max = 90.f ;
		:geospatial_lat_min = -90.f ;
		:geospatial_lat_resolution = "750 meters" ;
		:geospatial_lon_max = 180.f ;
		:geospatial_lon_min = -180.f ;
		:geospatial_lon_resolution = "750 meters" ;
		:id = "7c38eaa1-7e82-49dc-a00d-96fc30f77f4d" ;
		:geospatial_bounds = "POLYGON((92.3739319 -62.2583618, 17.40835 -73.4811554, 20.670002 -68.7148819, 84.2927856 -59.1303825, 92.3739319 -62.2583618))" ;
		:day_night_data_flag = "night" ;
		:start_orbit_number = 34108 ;
		:end_orbit_number = 34108 ;
		:ascend_descend_data_flag = 0 ;
		:geospatial_first_scanline_first_fov_lat = -62.25836f ;
		:geospatial_first_scanline_last_fov_lat = -59.13038f ;
		:geospatial_last_scanline_first_fov_lat = -73.48116f ;
		:geospatial_last_scanline_last_fov_lat = -68.71488f ;
		:geospatial_first_scanline_first_fov_lon = 92.37393f ;
		:geospatial_first_scanline_last_fov_lon = 84.29279f ;
		:geospatial_last_scanline_first_fov_lon = 17.40835f ;
		:geospatial_last_scanline_last_fov_lon = 20.67f ;
		:NCO = "netCDF Operators version 5.0.6 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco)" ;
data:

 IceConc =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, 67.32343, 84.27617, 69.62304, 58.03904, _, 
    75.2986, _, 93.43942, 89.14372, 90.32429,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, 69.33148, _, _, _, _, _, 92.32764, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 100, 100, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, 77.16252, _, 89.43716, _, 
    96.34447, 100, 100,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, 93.09033, _, 68.65797, 72.14285, 72.15576, _, _, _, _, _, 
    93.74178, _, 100, 100, 100,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 95.81432, _, _, _, 
    _, _, _, _, _, _, _, 83.46582, _, _, 70.99985, _, _, _, _, _, _, _, 
    90.44588, _, 100, 100,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 100, _, _, 
    _, _, 100, 100, _, _, _, _, _, _, _, _, _, _, _, _, 98.98752, 100, _, _, 
    100,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 100,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 87.24126, _, 100, _, 
    _, _, _, _, _, _, _, 88.74048, 91.04077, _, 73.66028, 77.14046, 72.86072, 
    _, 96.87101, _, 65.08202, _, 89.43575, _, 100, 100, 100,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, 69.14838, 74.81149, _, _, _, _, _, _, 92.22154, _, 
    100, 100, 100,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 100, _, _, 
    _, _, 100, _, _, _, _, _, _, _, _, _, _, _, _, _, 99.45397, _, _, 100, 100,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 100, _, _, 
    100, _, _, 100, 100, 90.56665, _, _, _, _, _, 87.64484, _, _, 91.27245, 
    _, 100, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    100, 100, _, _, _, 95.01587, _, 98.09937, 89.29044, _, _, _, 87.08566, 
    96.69353, 94.27303, _, _, 100, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 100, _, 
    _, _, _, 100, 98.30614, 94.49585, _, 95.56421, _, _, 91.44451, 94.2695, 
    93.61901, _, _, _, _, 100, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    100, 100, _, _, 100, _, _, 97.12012, _, _, _, _, 96.67687, _, 91.58325, 
    _, _, _, _, _, _ ;

 IceMap =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 2, 2, 0, 2, 0, 2, 2, 2,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 2, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 2, 0, 2, 2, 2,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 2, 0, 2, 2, 2, 0, 0, 0, 0, 0, 2, 0, 2, 2, 2,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 2, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 2, 0, 2, 2,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 
    0, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 0, 0, 2,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 2, 0, 0, 0, 0, 
    0, 0, 0, 0, 2, 2, 0, 2, 2, 2, 0, 2, 0, 2, 0, 2, 0, 2, 2, 2,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 2, 2, 0, 0, 0, 0, 0, 0, 2, 0, 2, 2, 2,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 
    0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 2, 2,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 2, 
    0, 0, 2, 2, 2, 0, 0, 0, 0, 0, 2, 0, 0, 2, 0, 2, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 
    2, 0, 0, 0, 2, 0, 2, 2, 0, 0, 0, 2, 2, 2, 0, 0, 2, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 
    0, 0, 2, 2, 2, 0, 2, 0, 0, 2, 2, 2, 0, 0, 0, 0, 2, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 
    2, 0, 0, 2, 0, 0, 2, 0, 0, 0, 0, 2, 0, 2, 0, 0, 0, 0, 0, 0 ;

 IceRetrPct = 92.00418 ;

 IceSrfTemp =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, 262.912, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, 262.748, 260.5441, 262.449, 263.9549, 
    _, 261.7112, _, 259.3529, 259.9113, 259.7578,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, 262.4869, _, _, _, _, _, 259.4974, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 258.0082, 258.4478, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, 261.4689, _, 259.8732, _, 
    258.9752, 258.0523, 257.7929,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, 259.8637, _, 262.5745, 262.1214, 262.1198, _, _, _, _, _, 
    259.3136, _, 258.0438, 257.6424, 257.6123,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 260.4814, _, _, _, 
    _, _, _, _, _, _, _, 261.0668, _, _, 262.27, _, _, _, _, _, _, _, 
    259.742, _, 257.781, 257.7041,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 259.4695, _, 
    _, _, _, 258.8402, 258.6626, _, _, _, _, _, _, _, _, _, _, _, _, 
    258.6316, 258.2289, _, _, 257.6414,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 257.6414,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 261.4673, _, 
    259.9039, _, _, _, _, _, _, _, _, 260.4074, 260.1199, _, 261.9242, 
    261.4717, 262.0281, _, 258.9068, _, 263.0393, _, 259.8734, _, 258.0083, 
    257.6029, 257.8393,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, 262.5107, 261.7745, _, _, _, _, _, _, 259.5112, _, 
    257.9245, 257.633, 257.3847,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 259.6055, _, 
    _, _, _, 258.671, _, _, _, _, _, _, _, _, _, _, _, _, _, 258.571, _, _, 
    257.6851, 257.6045,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 259.8718, _, 
    _, 259.1182, _, _, 259.2526, 259.4372, 260.1792, _, _, _, _, _, 260.1062, 
    _, _, 259.6346, _, 258.4996, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    259.1245, 259.1255, _, _, _, 259.623, _, 259.2376, 259.8922, _, _, _, 
    260.1789, 258.9298, 259.2445, _, _, 258.3249, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 259.6207, 
    _, _, _, _, 259.3116, 260.1948, 259.688, _, 259.5545, _, _, 259.6122, 
    259.245, 259.3295, _, _, _, _, 258.3306, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    259.3393, 259.3635, _, _, 259.6414, _, _, 259.36, _, _, _, _, 258.932, _, 
    259.5942, _, _, _, _, _, _ ;

 IceTermntPct = 96.45524 ;

 Latitude =
  -62.26201, -62.28693, -62.31173, -62.33637, -62.36088, -62.38528, 
    -62.40954, -62.43367, -62.45765, -62.48153, -62.50529, -62.52892, 
    -62.55244, -62.57583, -62.59911, -62.62225, -62.64531, -62.66823, 
    -62.69104, -62.71375, -62.73633, -62.7588, -62.78117, -62.80342, 
    -62.82558, -62.84762, -62.86955, -62.89139, -62.91312, -62.93473, 
    -62.95624, -62.97764, -62.99895, -63.02018, -63.04131, -63.06235, 
    -63.08331, -63.10412, -63.12487, -63.1455, -63.16606, -63.1865, 
    -63.20688, -63.22714, -63.24732,
  -62.24429, -62.26923, -62.29401, -62.31867, -62.34322, -62.36762, -62.3919, 
    -62.41604, -62.44005, -62.46393, -62.48772, -62.51137, -62.53489, 
    -62.5583, -62.5816, -62.60479, -62.62783, -62.65078, -62.6736, -62.69632, 
    -62.71892, -62.7414, -62.76378, -62.78606, -62.80823, -62.83027, 
    -62.85222, -62.87408, -62.89582, -62.91745, -62.93898, -62.96041, 
    -62.98171, -63.00295, -63.02411, -63.04518, -63.06613, -63.08697, 
    -63.10772, -63.12837, -63.14893, -63.1694, -63.18978, -63.21006, -63.23025,
  -62.22651, -62.25145, -62.27627, -62.30095, -62.32549, -62.34993, -62.3742, 
    -62.39836, -62.42241, -62.44631, -62.47009, -62.49377, -62.51731, 
    -62.54074, -62.56406, -62.58723, -62.61031, -62.63326, -62.65611, 
    -62.67884, -62.70145, -62.72396, -62.74635, -62.76864, -62.79083, 
    -62.81289, -62.83486, -62.85672, -62.87847, -62.90014, -62.92169, 
    -62.94311, -62.96445, -62.98568, -63.00685, -63.02795, -63.04889, 
    -63.06976, -63.09053, -63.11119, -63.13177, -63.15226, -63.17266, 
    -63.19294, -63.21315,
  -62.20868, -62.23362, -62.25846, -62.28316, -62.30772, -62.33216, 
    -62.35647, -62.38065, -62.40471, -62.42862, -62.45242, -62.4761, 
    -62.49968, -62.52313, -62.54646, -62.56966, -62.59274, -62.6157, 
    -62.63857, -62.66131, -62.68395, -62.70645, -62.72887, -62.75117, 
    -62.77337, -62.79546, -62.81743, -62.83931, -62.86109, -62.88277, 
    -62.90434, -62.92577, -62.94712, -62.96838, -62.98954, -63.01065, 
    -63.03164, -63.05252, -63.07329, -63.09396, -63.11456, -63.13505, 
    -63.15548, -63.17579, -63.196,
  -62.19078, -62.21574, -62.2406, -62.2653, -62.28989, -62.31435, -62.33867, 
    -62.36287, -62.38693, -62.41087, -62.4347, -62.45842, -62.48199, 
    -62.50544, -62.52879, -62.55201, -62.57511, -62.5981, -62.62097, 
    -62.64373, -62.66639, -62.68891, -62.71133, -62.73365, -62.75586, 
    -62.77798, -62.79998, -62.82188, -62.84368, -62.86536, -62.88693, 
    -62.90839, -62.92974, -62.95101, -62.97221, -62.99332, -63.01432, 
    -63.03521, -63.05601, -63.0767, -63.09731, -63.11782, -63.13824, 
    -63.15857, -63.17879,
  -62.17282, -62.19782, -62.22268, -62.2474, -62.272, -62.29648, -62.32082, 
    -62.34503, -62.36912, -62.39308, -62.41693, -62.44065, -62.46425, 
    -62.48772, -62.51107, -62.5343, -62.55743, -62.58043, -62.60332, 
    -62.6261, -62.64875, -62.67131, -62.69375, -62.71609, -62.73832, 
    -62.76044, -62.78246, -62.80437, -62.8262, -62.8479, -62.86947, 
    -62.89095, -62.91233, -62.9336, -62.95482, -62.97595, -62.99697, 
    -63.01787, -63.03868, -63.05939, -63.08001, -63.10055, -63.12098, 
    -63.14132, -63.16157,
  -62.15481, -62.17982, -62.20471, -62.22945, -62.25407, -62.27857, 
    -62.30292, -62.32715, -62.35126, -62.37523, -62.39909, -62.42284, 
    -62.44645, -62.46994, -62.4933, -62.51656, -62.5397, -62.56272, 
    -62.58563, -62.60842, -62.6311, -62.65367, -62.67613, -62.69849, 
    -62.72072, -62.74287, -62.76492, -62.78683, -62.80865, -62.83037, 
    -62.85198, -62.87346, -62.89486, -62.91616, -62.93738, -62.95853, 
    -62.97956, -63.00048, -63.02131, -63.04203, -63.06266, -63.08321, 
    -63.10367, -63.12402, -63.14428,
  -62.13674, -62.16177, -62.18667, -62.21144, -62.23608, -62.26059, 
    -62.28497, -62.30923, -62.33334, -62.35735, -62.38122, -62.40496, 
    -62.4286, -62.4521, -62.47549, -62.49877, -62.52193, -62.54496, 
    -62.56787, -62.59069, -62.61338, -62.63597, -62.65845, -62.68083, 
    -62.70309, -62.72525, -62.7473, -62.76923, -62.79108, -62.81281, 
    -62.83443, -62.85594, -62.87734, -62.89866, -62.9199, -62.94106, 
    -62.9621, -62.98305, -63.00388, -63.02463, -63.04528, -63.06583, 
    -63.0863, -63.10668, -63.12696,
  -62.20229, -62.22714, -62.25185, -62.27643, -62.3009, -62.32522, -62.34944, 
    -62.3735, -62.39744, -62.42127, -62.44497, -62.46856, -62.49202, 
    -62.51536, -62.53855, -62.56163, -62.58459, -62.60746, -62.63023, 
    -62.65292, -62.67546, -62.69792, -62.72024, -62.74243, -62.76454, 
    -62.78652, -62.80841, -62.83018, -62.85189, -62.87347, -62.89493, 
    -62.9163, -62.93758, -62.95876, -62.97982, -63.0008, -63.02162, 
    -63.04238, -63.06308, -63.08369, -63.1042, -63.1246, -63.14489, 
    -63.16511, -63.18526,
  -62.18449, -62.20935, -62.23409, -62.25868, -62.28314, -62.30751, 
    -62.33173, -62.35582, -62.37976, -62.4036, -62.42735, -62.45093, 
    -62.47441, -62.49775, -62.52097, -62.54407, -62.56704, -62.58994, 
    -62.61273, -62.6354, -62.65798, -62.68045, -62.70278, -62.725, -62.7471, 
    -62.76911, -62.79102, -62.81282, -62.83453, -62.85612, -62.8776, 
    -62.89899, -62.92028, -62.94146, -62.96255, -62.98352, -63.00439, 
    -63.02516, -63.04585, -63.06648, -63.08701, -63.10742, -63.12773, 
    -63.14795, -63.16812,
  -62.16662, -62.19151, -62.21626, -62.24088, -62.26535, -62.28973, 
    -62.31395, -62.33807, -62.36204, -62.38591, -62.40965, -62.43325, 
    -62.45674, -62.48012, -62.50335, -62.52645, -62.54944, -62.57235, 
    -62.59515, -62.61784, -62.64044, -62.66291, -62.68528, -62.7075, 
    -62.72963, -62.75167, -62.77359, -62.79539, -62.81711, -62.83872, 
    -62.86021, -62.88162, -62.90292, -62.92412, -62.94522, -62.96622, 
    -62.9871, -63.00787, -63.02859, -63.04924, -63.06976, -63.09018, 
    -63.11052, -63.13077, -63.15094,
  -62.1487, -62.17361, -62.19837, -62.22301, -62.2475, -62.27188, -62.29613, 
    -62.32028, -62.34426, -62.36814, -62.39189, -62.41552, -62.43902, 
    -62.46241, -62.48566, -62.50877, -62.5318, -62.55471, -62.57752, 
    -62.60024, -62.62286, -62.64535, -62.66772, -62.68998, -62.71213, 
    -62.73416, -62.75609, -62.77792, -62.79966, -62.82127, -62.84279, 
    -62.86421, -62.88552, -62.90673, -62.92785, -62.94887, -62.96976, 
    -62.99055, -63.01128, -63.03194, -63.05248, -63.07293, -63.09328, 
    -63.11353, -63.13371,
  -62.13073, -62.15564, -62.18042, -62.20507, -62.2296, -62.254, -62.27827, 
    -62.30242, -62.32643, -62.35032, -62.37409, -62.39773, -62.42126, 
    -62.44466, -62.46794, -62.49105, -62.51408, -62.53703, -62.55986, 
    -62.5826, -62.60523, -62.62773, -62.65012, -62.6724, -62.69455, 
    -62.71659, -62.73857, -62.7604, -62.78214, -62.80377, -62.82531, 
    -62.84675, -62.86807, -62.88932, -62.91044, -62.93147, -62.95238, 
    -62.97319, -62.99393, -63.01461, -63.03518, -63.05562, -63.07598, 
    -63.09626, -63.11648,
  -62.1127, -62.13765, -62.16243, -62.1871, -62.21166, -62.23609, -62.26037, 
    -62.28451, -62.30855, -62.33246, -62.35624, -62.3799, -62.40345, 
    -62.42686, -62.45015, -62.4733, -62.49633, -62.51929, -62.54214, 
    -62.56489, -62.58754, -62.61006, -62.63247, -62.65477, -62.67694, 
    -62.69901, -62.72098, -62.74283, -62.76459, -62.78625, -62.80779, 
    -62.82923, -62.85059, -62.87182, -62.89297, -62.91403, -62.93495, 
    -62.95576, -62.97654, -62.99721, -63.0178, -63.03827, -63.05866, 
    -63.07895, -63.09917,
  -62.0946, -62.11958, -62.1444, -62.16909, -62.19365, -62.21809, -62.24238, 
    -62.26656, -62.29061, -62.31452, -62.33832, -62.36201, -62.38557, 
    -62.40901, -62.43231, -62.45547, -62.47853, -62.5015, -62.52438, 
    -62.54714, -62.56981, -62.59236, -62.61476, -62.63708, -62.65927, 
    -62.68135, -62.70333, -62.7252, -62.74699, -62.76866, -62.79021, 
    -62.81168, -62.83305, -62.85431, -62.87547, -62.89653, -62.91748, 
    -62.93832, -62.95908, -62.97978, -63.00042, -63.0209, -63.04129, 
    -63.06158, -63.08181 ;

 Longitude =
  92.32836, 92.28934, 92.25043, 92.21167, 92.17303, 92.1345, 92.09612, 
    92.05786, 92.01971, 91.9817, 91.9438, 91.906, 91.86833, 91.83078, 
    91.79333, 91.75603, 91.7188, 91.68171, 91.64473, 91.60786, 91.57111, 
    91.53446, 91.4979, 91.46147, 91.42513, 91.38892, 91.35278, 91.31676, 
    91.28085, 91.24503, 91.20936, 91.17381, 91.13828, 91.10289, 91.06756, 
    91.0323, 90.99715, 90.96214, 90.92722, 90.8924, 90.85765, 90.82302, 
    90.78848, 90.75401, 90.71967,
  92.27644, 92.23746, 92.19865, 92.15996, 92.12137, 92.08293, 92.04461, 
    92.0064, 91.96834, 91.93037, 91.89256, 91.85484, 91.81721, 91.77973, 
    91.74236, 91.70508, 91.66795, 91.63094, 91.594, 91.5572, 91.52051, 
    91.48391, 91.44743, 91.41106, 91.37479, 91.33862, 91.30257, 91.26662, 
    91.23075, 91.19501, 91.15939, 91.12386, 91.08844, 91.05311, 91.01783, 
    90.98264, 90.94756, 90.9126, 90.87774, 90.84296, 90.80829, 90.77373, 
    90.73923, 90.70483, 90.67053,
  92.22459, 92.18573, 92.14696, 92.10833, 92.06983, 92.03144, 91.9932, 
    91.95507, 91.91708, 91.87918, 91.84142, 91.80374, 91.7662, 91.72879, 
    91.69146, 91.65427, 91.61721, 91.58024, 91.54339, 91.50665, 91.47001, 
    91.43347, 91.39709, 91.36076, 91.32457, 91.28845, 91.25244, 91.21656, 
    91.18079, 91.14509, 91.1095, 91.07404, 91.03868, 91.00343, 90.96821, 
    90.93306, 90.89806, 90.86316, 90.82837, 90.79366, 90.75903, 90.7245, 
    90.69007, 90.65573, 90.62152,
  92.17288, 92.13409, 92.09541, 92.05685, 92.01839, 91.98009, 91.9419, 
    91.90384, 91.8659, 91.82809, 91.79037, 91.75279, 91.71529, 91.67793, 
    91.64069, 91.60357, 91.56655, 91.52966, 91.49287, 91.45618, 91.41963, 
    91.38317, 91.34682, 91.31057, 91.27442, 91.23837, 91.20243, 91.16661, 
    91.13089, 91.09524, 91.05972, 91.02435, 90.98907, 90.95384, 90.91871, 
    90.88361, 90.84867, 90.81384, 90.77909, 90.74442, 90.70988, 90.67542, 
    90.64106, 90.60677, 90.5726,
  92.12129, 92.08257, 92.04397, 92.00547, 91.9671, 91.92885, 91.89072, 
    91.85273, 91.81487, 91.77711, 91.73946, 91.70191, 91.6645, 91.62721, 
    91.59003, 91.55297, 91.51604, 91.47919, 91.44247, 91.40585, 91.36934, 
    91.33295, 91.29668, 91.26048, 91.22441, 91.18842, 91.15255, 91.11676, 
    91.08108, 91.04552, 91.01008, 90.97475, 90.93951, 90.90437, 90.86929, 
    90.83427, 90.79936, 90.76458, 90.72989, 90.69531, 90.66081, 90.62642, 
    90.5921, 90.55789, 90.52377,
  92.06983, 92.03118, 91.99264, 91.95422, 91.91589, 91.87771, 91.83965, 
    91.80173, 91.76392, 91.72619, 91.68861, 91.65117, 91.61382, 91.57659, 
    91.53949, 91.5025, 91.46561, 91.42886, 91.39217, 91.35561, 91.31918, 
    91.28284, 91.24663, 91.21049, 91.17448, 91.13857, 91.10273, 91.06703, 
    91.03141, 90.9959, 90.96053, 90.92525, 90.89008, 90.855, 90.81996, 
    90.785, 90.75018, 90.71545, 90.68082, 90.64629, 90.61185, 90.57751, 
    90.54325, 90.50909, 90.47505,
  92.01849, 91.97987, 91.94141, 91.90305, 91.8648, 91.82668, 91.78869, 
    91.75083, 91.71306, 91.67544, 91.63794, 91.60052, 91.56325, 91.52608, 
    91.48905, 91.45212, 91.41531, 91.37858, 91.34199, 91.30551, 91.26913, 
    91.23284, 91.19669, 91.16062, 91.12466, 91.08879, 91.05303, 91.01737, 
    90.98183, 90.9464, 90.91106, 90.87588, 90.84076, 90.80573, 90.77076, 
    90.73586, 90.70107, 90.66644, 90.63184, 90.59737, 90.56301, 90.52871, 
    90.49451, 90.46043, 90.42643,
  91.96724, 91.92871, 91.8903, 91.85201, 91.81382, 91.77579, 91.73785, 
    91.70002, 91.66235, 91.62477, 91.58734, 91.55, 91.51279, 91.47569, 
    91.4387, 91.40185, 91.36508, 91.32845, 91.29192, 91.25548, 91.21917, 
    91.18296, 91.14687, 91.11082, 91.07494, 91.03915, 91.00345, 90.96786, 
    90.93236, 90.897, 90.86172, 90.82659, 90.79153, 90.75655, 90.72166, 
    90.68684, 90.6521, 90.6175, 90.583, 90.54856, 90.51425, 90.48003, 
    90.44591, 90.41185, 90.3779,
  92.14404, 92.10492, 92.06598, 92.02713, 91.98841, 91.94981, 91.91131, 
    91.87297, 91.83474, 91.79664, 91.75866, 91.72073, 91.68298, 91.64534, 
    91.60785, 91.5705, 91.53324, 91.49606, 91.45898, 91.42199, 91.3851, 
    91.34834, 91.31168, 91.27516, 91.23875, 91.20244, 91.16624, 91.13013, 
    91.0941, 91.05822, 91.02245, 90.98676, 90.95116, 90.91568, 90.88029, 
    90.84501, 90.80988, 90.77483, 90.73982, 90.70487, 90.67006, 90.63535, 
    90.60075, 90.56625, 90.5318,
  92.09234, 92.05331, 92.0144, 91.97564, 91.93698, 91.89843, 91.86002, 
    91.82175, 91.78358, 91.74553, 91.70758, 91.66977, 91.63207, 91.59453, 
    91.5571, 91.51981, 91.48261, 91.44552, 91.40848, 91.37154, 91.33472, 
    91.29803, 91.26144, 91.22499, 91.18864, 91.15239, 91.11625, 91.08018, 
    91.04424, 91.00842, 90.97269, 90.93704, 90.90154, 90.8661, 90.83077, 
    90.79557, 90.76048, 90.7255, 90.69056, 90.65569, 90.62093, 90.58629, 
    90.55173, 90.5173, 90.4829,
  92.04076, 92.00178, 91.96294, 91.92425, 91.88567, 91.8472, 91.80884, 
    91.77063, 91.73253, 91.69452, 91.65667, 91.61892, 91.58129, 91.54379, 
    91.50644, 91.46921, 91.4321, 91.39506, 91.35809, 91.32122, 91.28448, 
    91.24783, 91.2113, 91.17491, 91.13863, 91.10241, 91.06633, 91.03037, 
    90.99448, 90.9587, 90.92306, 90.88749, 90.85201, 90.81665, 90.78139, 
    90.74622, 90.71122, 90.67628, 90.64142, 90.60658, 90.57188, 90.53731, 
    90.50283, 90.46841, 90.43409,
  91.98926, 91.95037, 91.9116, 91.87297, 91.83447, 91.79605, 91.75777, 
    91.71959, 91.68156, 91.64364, 91.60586, 91.56818, 91.53062, 91.49319, 
    91.45589, 91.41873, 91.38167, 91.3447, 91.30782, 91.271, 91.23429, 
    91.19772, 91.16128, 91.12493, 91.08869, 91.05257, 91.01655, 90.98064, 
    90.94482, 90.90911, 90.8735, 90.83801, 90.8026, 90.7673, 90.73212, 
    90.697, 90.66203, 90.62717, 90.59236, 90.55759, 90.52296, 90.48843, 
    90.45401, 90.41969, 90.3854,
  91.93791, 91.89908, 91.8604, 91.82183, 91.78336, 91.74503, 91.70679, 
    91.66869, 91.63074, 91.59288, 91.55516, 91.51756, 91.48006, 91.4427, 
    91.40546, 91.36836, 91.33136, 91.29446, 91.25762, 91.22089, 91.18424, 
    91.14773, 91.11131, 91.07504, 91.03889, 91.00284, 90.96686, 90.93102, 
    90.89526, 90.85963, 90.82409, 90.78862, 90.75327, 90.71805, 90.68291, 
    90.64787, 90.61298, 90.57815, 90.5434, 90.5087, 90.47413, 90.43966, 
    90.40529, 90.37099, 90.33678,
  91.88667, 91.84789, 91.80927, 91.77076, 91.73237, 91.69408, 91.65593, 
    91.61791, 91.58001, 91.54224, 91.50457, 91.46703, 91.42961, 91.39231, 
    91.35513, 91.3181, 91.28117, 91.24432, 91.20754, 91.17088, 91.13429, 
    91.09781, 91.06149, 91.02528, 90.98918, 90.95319, 90.9173, 90.88151, 
    90.84582, 90.81021, 90.77474, 90.73937, 90.70409, 90.66892, 90.63383, 
    90.59882, 90.56401, 90.52924, 90.49453, 90.45992, 90.42538, 90.39097, 
    90.35665, 90.32244, 90.28828,
  91.83555, 91.79684, 91.75826, 91.71982, 91.6815, 91.64329, 91.60519, 
    91.56725, 91.52942, 91.49169, 91.45412, 91.41662, 91.37926, 91.34202, 
    91.30491, 91.26795, 91.23109, 91.19429, 91.15759, 91.12096, 91.08443, 
    91.04803, 91.01178, 90.97562, 90.9396, 90.90366, 90.86784, 90.83211, 
    90.79646, 90.76093, 90.72552, 90.69021, 90.65498, 90.61985, 90.58482, 
    90.5499, 90.51514, 90.48046, 90.44579, 90.41122, 90.37672, 90.34238, 
    90.30814, 90.27399, 90.23987 ;

 MaxIceConc = 100 ;

 MeanIceConc = 96.61342 ;

 MinIceConc = 7.335297 ;

 NumOfQACategories = 4 ;

 QCFlags =
  -16958209, -16958209, -16958209, -16958209, -16958209, -16958209, 
    -16958209, -16958209, -16958209, -16958209, -16958209, -16958209, 
    -16958209, -16958209, -18006798, -16958217, -16958209, -16958209, 
    -16958209, -16958209, -16958209, -16958209, -16958209, -16958209, 
    -16958209, -16958209, -16958209, -16958209, -16958209, -16958209, 
    -16958209, -16958209, -16958209, -16958209, -16958209, -22201095, 
    -22201104, -22201095, -22201104, -16958217, -22201095, -16958209, 
    -22201104, -22201104, -22201104,
  -16958209, -16958209, -16958209, -16958209, -16958209, -16958209, 
    -16958209, -16958209, -16958209, -16958209, -16958209, -16958209, 
    -16958209, -16958209, -16958209, -16958209, -16958209, -16958209, 
    -16958209, -16958209, -16958209, -16958209, -16958209, -16958209, 
    -16958209, -16958209, -16958209, -16958209, -16958209, -16958209, 
    -16958209, -16958209, -16958209, -16958209, -16958209, -16958217, 
    -16958209, -22201095, -16958209, -16958209, -16958209, -16958209, 
    -16958217, -22201095, -16958217,
  -16958209, -16958209, -16958209, -16958209, -16958209, -16958209, 
    -16958209, -16958209, -16958209, -16958209, -16958209, -16958209, 
    -16958209, -16958209, -16958209, -16958209, -16958209, -16958209, 
    -16958209, -16958209, -16958209, -16958209, -16958209, -16958209, 
    -16958209, -16958209, -16958209, -16958209, -16958209, -16958209, 
    -16958209, -16958209, -16958209, -16958209, -16958209, -16958209, 
    -16958217, -16958217, -16958217, -16958209, -16958217, -16958217, 
    -22201104, -22201095, -16958217,
  -16958209, -16958209, -16958209, -16958209, -16958209, -16958209, 
    -16958209, -16958209, -16958209, -16958209, -16958209, -16958209, 
    -16958209, -16958209, -16958209, -16958209, -16958209, -16958209, 
    -16958209, -16958209, -16958209, -16958209, -16958209, -16958209, 
    -16958209, -16958209, -16958209, -16958209, -16958209, -16958209, 
    -16958217, -16958209, -16958209, -16958209, -16958209, -16958217, 
    -16958209, -16958209, -22201095, -16958209, -22201104, -16958217, 
    -22201095, -22201095, -22201095,
  -16958209, -16958209, -16958209, -16958209, -16958209, -16958209, 
    -16958209, -16958209, -16958209, -16958209, -16958209, -16958209, 
    -16958209, -16958209, -16958209, -16958209, -16958209, -16958209, 
    -16958209, -16958209, -16958209, -16958209, -16958209, -16958209, 
    -16958209, -16958209, -16958209, -16958209, -16958209, -16958217, 
    -22201095, -16958217, -22201095, -22201104, -22201095, -16958217, 
    -16958217, -16958209, -16958209, -16958209, -22201095, -16958217, 
    -22201095, -22201104, -22201104,
  -16958209, -16958209, -16958209, -16958209, -16958209, -16958209, 
    -16958209, -16958209, -16958209, -16958209, -16958209, -16958209, 
    -16958209, -16958209, -16958209, -16958209, -16958209, -16958209, 
    -16958209, -22201095, -16958209, -16958209, -16958209, -16958209, 
    -16958209, -16958209, -16958209, -16958209, -16958209, -16958209, 
    -22201095, -16958209, -16958217, -22201095, -16958209, -16958217, 
    -16958209, -16958209, -16958217, -16958209, -16958217, -22201095, 
    -16958209, -22201104, -22201104,
  -16958209, -16958209, -16958209, -16958209, -16958209, -16958209, 
    -16958209, -16958209, -16958209, -16958209, -16958209, -16958209, 
    -16958209, -16958209, -16958209, -16958209, -16958209, -16958209, 
    -16958209, -16958209, -16958217, -22201095, -16958217, -16958209, 
    -16958209, -16958217, -22201095, -22201095, -16958209, -16958209, 
    -16958217, -16958217, -16958209, -16958209, -16958209, -16958209, 
    -16958209, -16958217, -16958217, -16958217, -22201095, -22201095, 
    -16958209, -16958209, -22201104,
  -16958209, -16958209, -16958209, -16958209, -16958209, -16958209, 
    -16958209, -16958209, -16958209, -16958209, -16958209, -16958209, 
    -16958209, -16958209, -16958209, -16958209, -16958209, -16958209, 
    -16958209, -16958209, -16958209, -16958209, -16958209, -16958209, 
    -16958209, -16958209, -16958209, -16958209, -16958209, -16958217, 
    -16958217, -16958209, -16958209, -16958209, -16958209, -16958209, 
    -16958209, -16958209, -16958209, -16958209, -16958217, -16958209, 
    -16958209, -16958209, -22201095,
  -16958209, -16958209, -16958209, -16958209, -16958209, -16958209, 
    -16958209, -16958209, -16958209, -16958209, -16958209, -16958209, 
    -16958209, -16958209, -16958209, -16958209, -16958209, -16958209, 
    -22201095, -16958209, -22201095, -16958209, -16958209, -16958209, 
    -16958209, -16958209, -16958209, -16958209, -16958209, -22201104, 
    -22201104, -16958217, -22201104, -22201104, -22201095, -16958209, 
    -22201095, -16958209, -22201104, -16958209, -22201104, -16958217, 
    -22201104, -22201095, -22201104,
  -16958209, -16958209, -16958209, -16958209, -16958209, -16958209, 
    -16958209, -16958209, -16958209, -16958209, -16958209, -16958209, 
    -16958209, -16958209, -16958209, -16958209, -16958209, -16958209, 
    -16958209, -16958209, -16958209, -16958209, -16958209, -16958209, 
    -16958209, -16958209, -16958209, -16958209, -16958209, -16958209, 
    -16958209, -16958217, -22201095, -22201095, -16958217, -16958209, 
    -16958209, -16958209, -16958217, -16958209, -22201095, -16958217, 
    -22201095, -22201104, -22201104,
  -16958209, -16958209, -16958209, -16958209, -16958209, -16958209, 
    -16958209, -16958209, -16958209, -16958209, -16958209, -16958209, 
    -16958209, -16958209, -16958209, -16958209, -16958209, -16958217, 
    -16958217, -16958209, -16958217, -22201095, -16958209, -16958209, 
    -16958209, -16958209, -22201095, -16958209, -16958209, -16958217, 
    -16958217, -16958209, -16958209, -16958209, -16958209, -16958209, 
    -16958209, -16958209, -16958209, -16958209, -22201095, -16958217, 
    -16958209, -22201104, -22201104,
  -16958209, -16958209, -16958209, -16958209, -16958209, -16958209, 
    -16958209, -16958209, -16958209, -16958209, -16958209, -16958209, 
    -16958209, -16958209, -16958209, -16958217, -16958217, -16958209, 
    -16958209, -16958209, -16958209, -22201095, -16958217, -16958217, 
    -22201095, -16958217, -16958209, -22201095, -22201095, -22201095, 
    -16958217, -16958217, -16958217, -16958209, -16958209, -22201095, 
    -16958209, -16958217, -22201104, -16958217, -22201095, -16958209, 
    -16958209, -16958209, -16958217,
  -16958209, -16958209, -16958209, -16958209, -16958209, -16958209, 
    -16958209, -16958209, -16958209, -16958209, -16958209, -16958209, 
    -16958209, -16958209, -16958217, -16958217, -16958217, -16958209, 
    -16958209, -16958209, -16958209, -16958209, -16958217, -16958217, 
    -22201095, -22201095, -16958217, -16958217, -16958217, -22201095, 
    -16958217, -22201095, -22201095, -16958209, -16958217, -16958209, 
    -22201095, -22201095, -22201104, -16958217, -16958217, -22201095, 
    -16958217, -16958209, -16958209,
  -16958209, -16958209, -16958209, -16958209, -16958209, -16958209, 
    -16958209, -16958209, -16958209, -16958209, -16958209, -16958209, 
    -16958209, -16958217, -16958209, -16958217, -16958217, -16958209, 
    -16958209, -16958209, -16958209, -16958209, -22201095, -16958217, 
    -16958217, -16958209, -16958217, -22201095, -22201095, -22201095, 
    -16958217, -22201104, -16958217, -16958217, -22201104, -22201095, 
    -22201104, -16958217, -16958209, -16958217, -16958209, -22201095, 
    -16958217, -16958209, -16958209,
  -16958209, -16958209, -16958209, -16958209, -16958209, -16958209, 
    -16958209, -16958209, -16958209, -16958209, -16958209, -16958209, 
    -16958209, -16958217, -16958217, -16958217, -16958217, -16958209, 
    -16958209, -16958209, -16958209, -16958209, -16958209, -16958217, 
    -22201095, -22201095, -16958217, -16958217, -22201095, -16958217, 
    -16958217, -22201095, -16958217, -16958217, -16958217, -16958217, 
    -22201095, -16958217, -22201095, -16958209, -16958217, -16958209, 
    -16958217, -16958209, -16958209 ;

 STDIceConc = 6.231885 ;

 SearchWindowSize = 50 ;

 StartColumn = 1 ;

 StartRow = 1 ;

 SummaryQC_Ice_Concentration =
  3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 2, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 
    3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 1, 0, 1, 0, 3, 1, 3, 0, 0, 0,
  3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 
    3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 1, 3, 3, 3, 3, 3, 1, 3,
  3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 
    3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 0, 1, 3,
  3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 
    3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 1, 3, 0, 3, 1, 1, 1,
  3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 
    3, 3, 3, 3, 3, 1, 3, 1, 0, 1, 3, 3, 3, 3, 3, 1, 3, 1, 0, 0,
  3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 1, 3, 3, 3, 3, 3, 
    3, 3, 3, 3, 3, 1, 3, 3, 1, 3, 3, 3, 3, 3, 3, 3, 1, 3, 0, 0,
  3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 1, 3, 3, 3, 
    3, 1, 1, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 1, 1, 3, 3, 0,
  3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 
    3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 1,
  3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 1, 3, 1, 3, 3, 3, 3, 
    3, 3, 3, 3, 0, 0, 3, 0, 0, 1, 3, 1, 3, 0, 3, 0, 3, 0, 1, 0,
  3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 
    3, 3, 3, 3, 3, 3, 3, 1, 1, 3, 3, 3, 3, 3, 3, 1, 3, 1, 0, 0,
  3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 1, 3, 3, 3, 
    3, 1, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 1, 3, 3, 0, 0,
  3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 1, 3, 3, 1, 
    3, 3, 1, 1, 1, 3, 3, 3, 3, 3, 1, 3, 3, 0, 3, 1, 3, 3, 3, 3,
  3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 1, 
    1, 3, 3, 3, 1, 3, 1, 1, 3, 3, 3, 1, 1, 0, 3, 3, 1, 3, 3, 3,
  3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 1, 3, 3, 
    3, 3, 1, 1, 1, 3, 0, 3, 3, 0, 1, 0, 3, 3, 3, 3, 1, 3, 3, 3,
  3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 1, 
    1, 3, 3, 1, 3, 3, 1, 3, 3, 3, 3, 1, 3, 1, 3, 3, 3, 3, 3, 3 ;

 TotDaytimePixs = _ ;

 TotIceRetrvls = 87116 ;

 TotIceTermnt = 2370484 ;

 TotNighttimePixs = 87116 ;

 TotWaterPixs = 94687 ;

 Tot_QA_BadData = 2362913 ;

 Tot_QA_Nonretrievable = 7571 ;

 Tot_QA_Normal = 37020 ;

 Tot_QA_Uncertain = 50096 ;

 cloud_mask_granule_level_quality_flag = 0 ;

 quality_information = 255 ;
}
