netcdf rads_adt_3a_2018104.tmp {
dimensions:
	time = UNLIMITED ; // (11 currently)
variables:
	int adt_egm2008(time) ;
		adt_egm2008:_FillValue = 2147483647 ;
		adt_egm2008:long_name = "absolute dynamic topography (EGM2008)" ;
		adt_egm2008:standard_name = "absolute_dynamic_topography_egm2008" ;
		adt_egm2008:units = "m" ;
		adt_egm2008:scale_factor = 0.0001 ;
		adt_egm2008:coordinates = "lon lat" ;
	int adt_xgm2016(time) ;
		adt_xgm2016:_FillValue = 2147483647 ;
		adt_xgm2016:long_name = "absolute dynamic topography (XGM2016)" ;
		adt_xgm2016:standard_name = "absolute_dynamic_topography_xgm2016" ;
		adt_xgm2016:units = "m" ;
		adt_xgm2016:scale_factor = 0.0001 ;
		adt_xgm2016:coordinates = "lon lat" ;
	int cycle(time) ;
		cycle:_FillValue = 2147483647 ;
		cycle:long_name = "cycle number" ;
		cycle:field = 9905s ;
	int lat(time) ;
		lat:_FillValue = 2147483647 ;
		lat:long_name = "latitude" ;
		lat:standard_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:scale_factor = 1.e-06 ;
		lat:field = 201s ;
		lat:comment = "Positive latitude is North latitude, negative latitude is South latitude" ;
	int lon(time) ;
		lon:_FillValue = 2147483647 ;
		lon:long_name = "longitude" ;
		lon:standard_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:scale_factor = 1.e-06 ;
		lon:field = 301s ;
		lon:comment = "East longitude relative to Greenwich meridian" ;
	int pass(time) ;
		pass:_FillValue = 2147483647 ;
		pass:long_name = "pass number" ;
		pass:field = 9906s ;
	short sla(time) ;
		sla:_FillValue = 32767s ;
		sla:long_name = "sea level anomaly" ;
		sla:standard_name = "sea_surface_height_above_sea_level" ;
		sla:units = "m" ;
		sla:quality_flag = "swh sig0 range_rms range_numval flags swh_rms sig0_rms" ;
		sla:scale_factor = 0.0001 ;
		sla:coordinates = "lon lat" ;
		sla:field = 0s ;
		sla:comment = "Sea level determined from satellite altitude - range - all altimetric corrections" ;
	double time_mjd(time) ;
		time_mjd:long_name = "Modified Julian Days" ;
		time_mjd:standard_name = "time" ;
		time_mjd:units = "days since 1858-11-17 00:00:00 UTC" ;
		time_mjd:field = 105s ;
		time_mjd:comment = "UTC time of measurement expressed in Modified Julian Days" ;

// global attributes:
		:Conventions = "CF-1.7" ;
		:title = "RADS 4 pass file" ;
		:institution = "EUMETSAT / NOAA / TU Delft" ;
		:source = "radar altimeter" ;
		:references = "RADS Data Manual, Version 4.2 or later" ;
		:featureType = "trajectory" ;
		:ellipsoid = "TOPEX" ;
		:ellipsoid_axis = 6378136.3 ;
		:ellipsoid_flattening = 0.00335281317789691 ;
		:filename = "rads_adt_3a_2018104.nc" ;
		:mission_name = "SNTNL-3A" ;
		:mission_phase = "a" ;
		:log01 = "2019-01-11 | rads2nc --ymd=180414000000,180415000000 -C1,1000 -S3a -Vadt_egm2008,adt_xgm2016,sla,time_mjd,lon,lat,cycle,pass -Xxgm2016 -Xadt.xml -o/ftp/rads/adt//2018/rads_adt_3a_2018104.nc: RAW data from" ;
		:history = "Fri Jan 26 15:44:21 2024: ncks -d time,0,10 /scratch1/NCEPDEV/stmp4/Shastri.Paturi/forAndrew/gdas.20180414/00/adt/rads_adt_3a_2018104.nc rads_adt_3a_2018104.tmp.nc\n",
			"2019-01-11 12:29:34 : rads2nc --ymd=180414000000,180415000000 -C1,1000 -S3a -Vadt_egm2008,adt_xgm2016,sla,time_mjd,lon,lat,cycle,pass -Xxgm2016 -Xadt.xml -o/ftp/rads/adt//2018/rads_adt_3a_2018104.nc" ;
		:NCO = "netCDF Operators version 5.0.6 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco)" ;
data:

 adt_egm2008 = -10834, -11080, -11752, -12215, -12322, -12631, -12835, 
    -13106, -13520, -13476, -13197 ;

 adt_xgm2016 = -11476, -10955, -12265, -13723, -13874, -13752, -13406, 
    -13319, -13383, -13127, -12743 ;

 cycle = 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30 ;

 lat = -68340968, -68286987, -68232981, -68178950, -68124894, -68070813, 
    -68016708, -67962578, -67908424, -67854245, -67800043 ;

 lon = -8586260, -8654949, -8723334, -8791417, -8859200, -8926685, -8993875, 
    -9060771, -9127375, -9193690, -9259717 ;

 pass = 175, 175, 175, 175, 175, 175, 175, 175, 175, 175, 175 ;

 sla = 347, 463, 323, 207, 153, 107, 174, -96, -252, -8, 527 ;

 time_mjd = 58222.0026388889, 58222.002650463, 58222.002662037, 
    58222.0026736111, 58222.0026851852, 58222.0026967593, 58222.0027083333, 
    58222.0027199074, 58222.0027314815, 58222.0027430556, 58222.0027546296 ;
}
