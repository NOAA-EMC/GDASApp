netcdf rads_adt_sa_2018105.tmp {
dimensions:
	time = UNLIMITED ; // (11 currently)
variables:
	int adt_egm2008(time) ;
		adt_egm2008:_FillValue = 2147483647 ;
		adt_egm2008:long_name = "absolute dynamic topography (EGM2008)" ;
		adt_egm2008:standard_name = "absolute_dynamic_topography_egm2008" ;
		adt_egm2008:units = "m" ;
		adt_egm2008:scale_factor = 0.0001 ;
		adt_egm2008:coordinates = "lon lat" ;
	int adt_xgm2016(time) ;
		adt_xgm2016:_FillValue = 2147483647 ;
		adt_xgm2016:long_name = "absolute dynamic topography (XGM2016)" ;
		adt_xgm2016:standard_name = "absolute_dynamic_topography_xgm2016" ;
		adt_xgm2016:units = "m" ;
		adt_xgm2016:scale_factor = 0.0001 ;
		adt_xgm2016:coordinates = "lon lat" ;
	int cycle(time) ;
		cycle:_FillValue = 2147483647 ;
		cycle:long_name = "cycle number" ;
		cycle:field = 9905s ;
	int lat(time) ;
		lat:_FillValue = 2147483647 ;
		lat:long_name = "latitude" ;
		lat:standard_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:scale_factor = 1.e-06 ;
		lat:field = 201s ;
		lat:comment = "Positive latitude is North latitude, negative latitude is South latitude" ;
	int lon(time) ;
		lon:_FillValue = 2147483647 ;
		lon:long_name = "longitude" ;
		lon:standard_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:scale_factor = 1.e-06 ;
		lon:field = 301s ;
		lon:comment = "East longitude relative to Greenwich meridian" ;
	int pass(time) ;
		pass:_FillValue = 2147483647 ;
		pass:long_name = "pass number" ;
		pass:field = 9906s ;
	short sla(time) ;
		sla:_FillValue = 32767s ;
		sla:long_name = "sea level anomaly" ;
		sla:standard_name = "sea_surface_height_above_sea_level" ;
		sla:units = "m" ;
		sla:quality_flag = "swh sig0 range_rms range_numval flags peakiness" ;
		sla:scale_factor = 0.0001 ;
		sla:coordinates = "lon lat" ;
		sla:field = 0s ;
		sla:comment = "Sea level determined from satellite altitude - range - all altimetric corrections" ;
	double time_mjd(time) ;
		time_mjd:long_name = "Modified Julian Days" ;
		time_mjd:standard_name = "time" ;
		time_mjd:units = "days since 1858-11-17 00:00:00 UTC" ;
		time_mjd:field = 105s ;
		time_mjd:comment = "UTC time of measurement expressed in Modified Julian Days" ;

// global attributes:
		:Conventions = "CF-1.7" ;
		:title = "RADS 4 pass file" ;
		:institution = "EUMETSAT / NOAA / TU Delft" ;
		:source = "radar altimeter" ;
		:references = "RADS Data Manual, Version 4.2 or later" ;
		:featureType = "trajectory" ;
		:ellipsoid = "TOPEX" ;
		:ellipsoid_axis = 6378136.3 ;
		:ellipsoid_flattening = 0.00335281317789691 ;
		:filename = "rads_adt_sa_2018105.nc" ;
		:mission_name = "SARAL" ;
		:mission_phase = "b" ;
		:log01 = "2019-01-11 | rads2nc --ymd=180415000000,180416000000 -C1,1000 -Ssa -Vadt_egm2008,adt_xgm2016,sla,time_mjd,lon,lat,cycle,pass -Xxgm2016 -Xadt.xml -o/ftp/rads/adt//2018/rads_adt_sa_2018105.nc: RAW data from" ;
		:history = "Fri Jan 26 15:41:52 2024: ncks -d time,0,10 /scratch1/NCEPDEV/stmp4/Shastri.Paturi/forAndrew/gdas.20180415/00/adt/rads_adt_sa_2018105.nc rads_adt_sa_2018105.tmp.nc\n",
			"2019-01-11 12:29:44 : rads2nc --ymd=180415000000,180416000000 -C1,1000 -Ssa -Vadt_egm2008,adt_xgm2016,sla,time_mjd,lon,lat,cycle,pass -Xxgm2016 -Xadt.xml -o/ftp/rads/adt//2018/rads_adt_sa_2018105.nc" ;
		:NCO = "netCDF Operators version 5.0.6 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco)" ;
data:

 adt_egm2008 = 4713, 4144, 4098, 4152, 3662, 3363, 4196, 4149, 4308, 3574, 
    3516 ;

 adt_xgm2016 = 5346, 5058, 5316, 5518, 5322, 5182, 5536, 4657, 3992, 2985, 
    3213 ;

 cycle = 54, 54, 54, 54, 54, 54, 54, 54, 54, 54, 54 ;

 lat = 41652607, 41591789, 41530967, 41470143, 41409315, 41348485, 41287651, 
    41226815, 41165976, 41105134, 41044289 ;

 lon = -124261530, -124282255, -124302949, -124323613, -124344246, 
    -124364849, -124385422, -124405964, -124426477, -124446960, -124467413 ;

 pass = 558, 558, 558, 558, 558, 558, 558, 558, 558, 558, 558 ;

 sla = 580, 59, -82, -382, -567, -779, 2, 2, 170, -774, -581 ;

 time_mjd = 58223.1157344669, 58223.1157464813, 58223.1157584958, 
    58223.1157705102, 58223.1157825246, 58223.1157945391, 58223.1158065535, 
    58223.115818568, 58223.1158305824, 58223.1158425969, 58223.1158546113 ;
}
