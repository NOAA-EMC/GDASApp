netcdf rads_adt_j2_2018104.tmp {
dimensions:
	time = UNLIMITED ; // (11 currently)
variables:
	int adt_egm2008(time) ;
		adt_egm2008:_FillValue = 2147483647 ;
		adt_egm2008:long_name = "absolute dynamic topography (EGM2008)" ;
		adt_egm2008:standard_name = "absolute_dynamic_topography_egm2008" ;
		adt_egm2008:units = "m" ;
		adt_egm2008:scale_factor = 0.0001 ;
		adt_egm2008:coordinates = "lon lat" ;
	int adt_xgm2016(time) ;
		adt_xgm2016:_FillValue = 2147483647 ;
		adt_xgm2016:long_name = "absolute dynamic topography (XGM2016)" ;
		adt_xgm2016:standard_name = "absolute_dynamic_topography_xgm2016" ;
		adt_xgm2016:units = "m" ;
		adt_xgm2016:scale_factor = 0.0001 ;
		adt_xgm2016:coordinates = "lon lat" ;
	int cycle(time) ;
		cycle:_FillValue = 2147483647 ;
		cycle:long_name = "cycle number" ;
		cycle:field = 9905s ;
	int lat(time) ;
		lat:_FillValue = 2147483647 ;
		lat:long_name = "latitude" ;
		lat:standard_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:scale_factor = 1.e-06 ;
		lat:field = 201s ;
		lat:comment = "Positive latitude is North latitude, negative latitude is South latitude" ;
	int lon(time) ;
		lon:_FillValue = 2147483647 ;
		lon:long_name = "longitude" ;
		lon:standard_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:scale_factor = 1.e-06 ;
		lon:field = 301s ;
		lon:comment = "East longitude relative to Greenwich meridian" ;
	int pass(time) ;
		pass:_FillValue = 2147483647 ;
		pass:long_name = "pass number" ;
		pass:field = 9906s ;
	short sla(time) ;
		sla:_FillValue = 32767s ;
		sla:long_name = "sea level anomaly" ;
		sla:standard_name = "sea_surface_height_above_sea_level" ;
		sla:units = "m" ;
		sla:quality_flag = "swh sig0 range_rms range_numval flags swh_rms sig0_rms attitude" ;
		sla:scale_factor = 0.0001 ;
		sla:coordinates = "lon lat" ;
		sla:field = 0s ;
		sla:comment = "Sea level determined from satellite altitude - range - all altimetric corrections" ;
	double time_mjd(time) ;
		time_mjd:long_name = "Modified Julian Days" ;
		time_mjd:standard_name = "time" ;
		time_mjd:units = "days since 1858-11-17 00:00:00 UTC" ;
		time_mjd:field = 105s ;
		time_mjd:comment = "UTC time of measurement expressed in Modified Julian Days" ;

// global attributes:
		:Conventions = "CF-1.7" ;
		:title = "RADS 4 pass file" ;
		:institution = "EUMETSAT / NOAA / TU Delft" ;
		:source = "radar altimeter" ;
		:references = "RADS Data Manual, Version 4.2 or later" ;
		:featureType = "trajectory" ;
		:ellipsoid = "TOPEX" ;
		:ellipsoid_axis = 6378136.3 ;
		:ellipsoid_flattening = 0.00335281317789691 ;
		:filename = "rads_adt_j2_2018104.nc" ;
		:mission_name = "JASON-2" ;
		:mission_phase = "c" ;
		:log01 = "2019-01-11 | rads2nc --ymd=180414000000,180415000000 -C1,1000 -Sj2 -Vadt_egm2008,adt_xgm2016,sla,time_mjd,lon,lat,cycle,pass -Xxgm2016 -Xadt.xml -o/ftp/rads/adt//2018/rads_adt_j2_2018104.nc: RAW data from" ;
		:history = "Fri Jan 26 15:44:21 2024: ncks -d time,0,10 /scratch1/NCEPDEV/stmp4/Shastri.Paturi/forAndrew/gdas.20180414/00/adt/rads_adt_j2_2018104.nc rads_adt_j2_2018104.tmp.nc\n",
			"2019-01-11 12:29:31 : rads2nc --ymd=180414000000,180415000000 -C1,1000 -Sj2 -Vadt_egm2008,adt_xgm2016,sla,time_mjd,lon,lat,cycle,pass -Xxgm2016 -Xadt.xml -o/ftp/rads/adt//2018/rads_adt_j2_2018104.nc" ;
		:NCO = "netCDF Operators version 5.0.6 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco)" ;
data:

 adt_egm2008 = 9986, 10036, 9510, 9672, 9964, 9707, 9823, 9672, 9731, 9720, 
    9506 ;

 adt_xgm2016 = 8982, 9545, 9435, 10130, 10467, 9827, 9687, 9405, 9201, 9110, 
    8949 ;

 cycle = 349, 349, 349, 349, 349, 349, 349, 349, 349, 349, 349 ;

 lat = 10287080, 10238060, 10189039, 10140015, 10090990, 10041963, 9992935, 
    9943904, 9894873, 9845839, 9796804 ;

 lon = -177073813, -177055552, -177037298, -177019051, -177000811, 
    -176982578, -176964351, -176946131, -176927918, -176909711, -176891511 ;

 pass = 82, 82, 82, 82, 82, 82, 82, 82, 82, 82, 82 ;

 sla = 702, 799, 347, 458, 860, 709, 845, 776, 808, 710, 658 ;

 time_mjd = 58222.0000087827, 58222.0000203326, 58222.0000318827, 
    58222.0000434327, 58222.0000549827, 58222.0000665327, 58222.0000780827, 
    58222.0000896326, 58222.0001011826, 58222.0001127326, 58222.0001242827 ;
}
