netcdf icec.nc {
dimensions:
	Location = 100 ;
	nvars = 1 ;
variables:
	int Location(Location) ;
		Location:suggested_chunk_dim = 100LL ;
	float nvars(nvars) ;
		nvars:suggested_chunk_dim = 100LL ;

// global attributes:
		string :_ioda_layout = "ObsGroup" ;
		:_ioda_layout_version = 0 ;
		:converter = "somthing.py" ;
		:nvars = 1 ;
		:date_time = 2018041512 ;
		:nlocs = 100 ;
		:nobs = 100 ;
		:history = "Wed May 12 11:02:49 2021: ncks -O -4 icec.nc icec.nc4" ;
		:NCO = "netCDF Operators version 4.7.9 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco)" ;
data:

 Location = 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0 ;

 nvars = 0 ;

group: MetaData {
  variables:
  	int64 dateTime(Location) ;
  		dateTime:_FillValue = -2208988800LL ;
  		string dateTime:units = "seconds since 1970-01-01T00:00:00Z" ;
  	float latitude(Location) ;
  		latitude:_FillValue = 9.96921e+36f ;
  	float longitude(Location) ;
  		longitude:_FillValue = 9.96921e+36f ;
  	string variable_names(nvars) ;
  		string variable_names:_FillValue = "" ;
  data:

   dateTime = 1523756403, 1523755138, 1523809850, 1523761241, 1523822234, 
      1523768790, 1523785038, 1523759437, 1523766482, 1523810666, 1523796805, 
      1523793968, 1523823489, 1523752584, 1523775969, 1523762155, 1523768587, 
      1523814065, 1523804452, 1523785153, 1523814803, 1523798982, 1523809343, 
      1523817342, 1523781349, 1523820098, 1523791041, 1523769787, 1523815706, 
      1523778971, 1523804767, 1523796237, 1523824707, 1523818565, 1523751405, 
      1523787456, 1523810909, 1523762957, 1523791035, 1523792510, 1523786864, 
      1523790617, 1523814394, 1523791642, 1523755808, 1523810550, 1523762563, 
      1523777575, 1523781304, 1523777512, 1523783413, 1523800295, 1523767606, 
      1523780294, 1523787500, 1523805171, 1523833527, 1523761005, 1523774017, 
      1523834116, 1523751669, 1523750758, 1523755978, 1523756554, 1523801484, 
      1523818162, 1523824621, 1523818222, 1523806101, 1523766245, 1523832461, 
      1523793475, 1523804854, 1523775300, 1523766009, 1523777548, 1523817482, 
      1523779036, 1523830924, 1523807451, 1523821977, 1523793607, 1523832064, 
      1523814637, 1523802742, 1523807362, 1523807507, 1523802980, 1523780526, 
      1523795959, 1523758548, 1523761287, 1523830764, 1523831286, 1523762363, 
      1523833304, 1523750667, 1523809587, 1523760587, 1523798073 ;

   latitude = -78.375, -77.375, -76.625, -76.125, -75.625, -75.125, -74.875, 
      -74.375, -74.125, -73.625, -73.375, -72.875, -72.625, -72.375, -72.125, 
      -71.875, -71.625, -71.375, -70.875, -70.625, -70.375, -70.125, -69.875, 
      -69.625, -69.375, -69.125, -68.625, -68.375, -68.125, -67.625, -66.875, 
      -66.375, -66.125, -65.625, -65.375, -64.875, -64.375, -63.125, 49.125, 
      52.625, 55.125, 57.125, 58.875, 60.375, 61.875, 63.125, 64.375, 65.625, 
      67.125, 67.875, 68.625, 69.375, 69.875, 70.375, 70.625, 71.125, 71.625, 
      72.125, 72.375, 72.875, 73.375, 73.875, 74.375, 74.875, 75.375, 75.875, 
      76.125, 76.375, 76.875, 77.125, 77.375, 77.625, 77.875, 78.125, 78.625, 
      78.875, 79.125, 79.375, 79.625, 79.875, 80.375, 80.625, 80.875, 81.125, 
      81.375, 81.625, 81.875, 82.125, 82.375, 82.875, 83.125, 83.375, 83.875, 
      84.125, 84.625, 84.875, 85.375, 85.625, 85.875, 86.125 ;

   longitude = 178.625, 185.875, 163.125, 184.625, 193.125, 184.375, 334.375, 
      224.125, 339.375, 221.875, 315.125, 180.125, 217.375, 242.625, 269.625, 
      284.125, 322.625, 337.375, 179.125, 195.625, 231.375, 243.125, 256.375, 
      285.875, 314.875, 353.125, 4.375, 73.125, 311.875, 315.375, 68.375, 
      76.625, 300.625, 83.875, 142.625, 92.375, 116.875, 309.875, 306.625, 
      145.875, 147.625, 143.625, 158.875, 159.375, 276.875, 297.125, 195.375, 
      181.375, 73.375, 336.625, 295.375, 56.625, 162.375, 55.625, 299.625, 
      238.125, 190.625, 49.625, 284.875, 339.625, 344.625, 263.375, 128.375, 
      21.625, 75.875, 32.625, 150.125, 277.625, 14.375, 34.375, 58.375, 
      93.875, 165.875, 254.125, 23.875, 46.125, 63.125, 101.125, 160.625, 
      294.875, 38.625, 80.875, 119.625, 153.125, 156.875, 182.375, 197.375, 
      271.375, 346.625, 24.125, 151.125, 318.875, 107.125, 176.375, 131.875, 
      187.375, 3.375, 144.875, 164.625, 251.625 ;

   variable_names = "sea_ice_area_fraction" ;
  } // group MetaData

group: ObsError {
  variables:
  	float seaIceFraction(Location) ;
  		seaIceFraction:_FillValue = 9.96921e+36f ;
  data:

   seaIceFraction = 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 
      0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 
      0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 
      0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 
      0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 
      0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 
      0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 0.1, 
      0.1, 0.1, 0.1, 0.1, 0.1 ;
  } // group ObsError

group: ObsValue {
  variables:
  	float seaIceFraction(Location) ;
  		seaIceFraction:_FillValue = 9.96921e+36f ;
  data:

   seaIceFraction = 0.66, 0.86, 0.72, 0.94, 0.92, 0.94, 0.7, 0.72, 0.65, 
      0.81, 0.89, 0.87, 0.59, 0.89, 0.81, 0.51, 0.88, 0.32, 0.76, 0.78, 0.4, 
      0.4, 0.74, 0.52, 0.81, 0.48, 0.35, 0.66, 0.83, 0.72, 0.62, 0.78, 0.86, 
      0.8, 0.35, 0.64, 0.25, 0.39, 0.28, 0.72, 0.25, 0.96, 0.21, 0.26, 
      0.9899999, 0.98, 0.67, 0.39, 0.97, 0.33, 0.98, 0.77, 0.9899999, 0.66, 
      0.9899999, 0.9899999, 0.9899999, 0.22, 0.74, 0.92, 0.65, 0.9899999, 
      0.9899999, 0.38, 0.9899999, 0.22, 0.98, 0.98, 0.3, 0.8, 0.85, 0.98, 
      0.96, 0.9899999, 0.84, 0.93, 0.9899999, 0.84, 0.98, 0.8, 0.95, 
      0.9899999, 0.9899999, 0.9899999, 0.9899999, 0.98, 0.9899999, 0.94, 
      0.9899999, 0.9899999, 0.9899999, 0.9899999, 0.9899999, 0.9899999, 
      0.9899999, 0.9899999, 0.98, 0.9899999, 0.9899999, 0.9899999 ;
  } // group ObsValue

group: PreQc {
  variables:
  	float seaIceFraction(Location) ;
  		seaIceFraction:_FillValue = 9.96921e+36f ;
  data:

   seaIceFraction = 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
      0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
      0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
      0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
      0, 0, 0, 0, 0, 0, 0, 0, 0 ;
  } // group PreQc
}
