netcdf sss_smos_2 {
dimensions:
	n_grid_points = 52 ;
variables:
	float A_card(n_grid_points) ;
		A_card:_FillValue = -999.f ;
	ubyte Coast_distance(n_grid_points) ;
		Coast_distance:_FillValue = 0UB ;
		Coast_distance:scale_factor = 20. ;
		Coast_distance:scale_offset = 0. ;
		string Coast_distance:_Unsigned = "true" ;
	uint Control_Flags_Acard(n_grid_points) ;
		Control_Flags_Acard:_FillValue = 0U ;
		Control_Flags_Acard:flag_masks = 2s, 4s, 8s, 16s, 32s, 64s, 128s, 256s, 512s, 1024s, 2048s, 4096s, 8192s, 16384s, -32768s, 0s, 0s, 0s, 0s, 0s, 0s, 0s, 0s, 0s, 0s, 0s, 0s, 0s, 0s ;
		Control_Flags_Acard:flag_values = 2s, 4s, 8s, 16s, 32s, 64s, 128s, 256s, 512s, 1024s, 2048s, 4096s, 8192s, 16384s, -32768s, 0s, 0s, 0s, 0s, 0s, 0s, 0s, 0s, 0s, 0s, 0s, 0s, 0s, 0s ;
		string Control_Flags_Acard:flag_meanings = "FG_CTRL_RANGE FG_CTRL_SIGMA FG_CTRL_CHI2 FG_CTRL_CHI2_P FG_CTRL_CONTAMINATED FG_CTRL_SUNGLINT FG_CTRL_MOONGLINT FG_CTRL_GAL_NOISE FG_CTRL_MIXED_SCENE FG_CTRL_REACH_MAXITER FG_CTRL_NUM_MEAS_MIN FG_CTRL_NUM_MEAS_LOW FG_CTRL_MANY_OUTLIERS FG_CTRL_MARQ FG_CTRL_ROUGHNESS FG_CTRL_FOAM FG_CTRL_ECMWF FG_CTRL_VALID FG_CTRL_NO_SURFACE FG_CTRL_RANGE_ACARD FG_CTRL_SIGMA_ACARD FG_CTRL_USED_FARATEC FG_CTRL_POOR_GEOPHYS FG_CTRL_POOR_RETRIEVAL FG_CTRL_SUSPECT_RFI FG_CTRL_RFI_PRONE_X FG_CTRL_RFI_PRONE_Y FG_CTRL_ADJUSTED_RA FG_CTRL_RETRIEV_FAIL" ;
		string Control_Flags_Acard:_Unsigned = "true" ;
	uint Control_Flags_anom(n_grid_points) ;
		Control_Flags_anom:_FillValue = 0U ;
		Control_Flags_anom:flag_masks = 2s, 4s, 8s, 16s, 32s, 64s, 128s, 256s, 512s, 1024s, 2048s, 4096s, 8192s, 16384s, -32768s, 0s, 0s, 0s, 0s, 0s, 0s, 0s, 0s, 0s, 0s, 0s, 0s, 0s, 0s ;
		Control_Flags_anom:flag_values = 2s, 4s, 8s, 16s, 32s, 64s, 128s, 256s, 512s, 1024s, 2048s, 4096s, 8192s, 16384s, -32768s, 0s, 0s, 0s, 0s, 0s, 0s, 0s, 0s, 0s, 0s, 0s, 0s, 0s, 0s ;
		string Control_Flags_anom:flag_meanings = "FG_CTRL_RANGE FG_CTRL_SIGMA FG_CTRL_CHI2 FG_CTRL_CHI2_P FG_CTRL_CONTAMINATED FG_CTRL_SUNGLINT FG_CTRL_MOONGLINT FG_CTRL_GAL_NOISE FG_CTRL_MIXED_SCENE FG_CTRL_REACH_MAXITER FG_CTRL_NUM_MEAS_MIN FG_CTRL_NUM_MEAS_LOW FG_CTRL_MANY_OUTLIERS FG_CTRL_MARQ FG_CTRL_ROUGHNESS FG_CTRL_FOAM FG_CTRL_ECMWF FG_CTRL_VALID FG_CTRL_NO_SURFACE FG_CTRL_RANGE_ACARD FG_CTRL_SIGMA_ACARD FG_CTRL_USED_FARATEC FG_CTRL_POOR_GEOPHYS FG_CTRL_POOR_RETRIEVAL FG_CTRL_SUSPECT_RFI FG_CTRL_RFI_PRONE_X FG_CTRL_RFI_PRONE_Y FG_CTRL_ADJUSTED_RA FG_CTRL_RETRIEV_FAIL" ;
		string Control_Flags_anom:_Unsigned = "true" ;
	uint Control_Flags_corr(n_grid_points) ;
		Control_Flags_corr:_FillValue = 0U ;
		Control_Flags_corr:flag_masks = 2s, 4s, 8s, 16s, 32s, 64s, 128s, 256s, 512s, 1024s, 2048s, 4096s, 8192s, 16384s, -32768s, 0s, 0s, 0s, 0s, 0s, 0s, 0s, 0s, 0s, 0s, 0s, 0s, 0s, 0s ;
		Control_Flags_corr:flag_values = 2s, 4s, 8s, 16s, 32s, 64s, 128s, 256s, 512s, 1024s, 2048s, 4096s, 8192s, 16384s, -32768s, 0s, 0s, 0s, 0s, 0s, 0s, 0s, 0s, 0s, 0s, 0s, 0s, 0s, 0s ;
		string Control_Flags_corr:flag_meanings = "FG_CTRL_RANGE FG_CTRL_SIGMA FG_CTRL_CHI2 FG_CTRL_CHI2_P FG_CTRL_CONTAMINATED FG_CTRL_SUNGLINT FG_CTRL_MOONGLINT FG_CTRL_GAL_NOISE FG_CTRL_MIXED_SCENE FG_CTRL_REACH_MAXITER FG_CTRL_NUM_MEAS_MIN FG_CTRL_NUM_MEAS_LOW FG_CTRL_MANY_OUTLIERS FG_CTRL_MARQ FG_CTRL_ROUGHNESS FG_CTRL_FOAM FG_CTRL_ECMWF FG_CTRL_VALID FG_CTRL_NO_SURFACE FG_CTRL_RANGE_ACARD FG_CTRL_SIGMA_ACARD FG_CTRL_USED_FARATEC FG_CTRL_POOR_GEOPHYS FG_CTRL_POOR_RETRIEVAL FG_CTRL_SUSPECT_RFI FG_CTRL_RFI_PRONE_X FG_CTRL_RFI_PRONE_Y FG_CTRL_ADJUSTED_RA FG_CTRL_RETRIEV_FAIL" ;
		string Control_Flags_corr:_Unsigned = "true" ;
	uint Control_Flags_uncorr(n_grid_points) ;
		Control_Flags_uncorr:_FillValue = 0U ;
		Control_Flags_uncorr:flag_masks = 2s, 4s, 8s, 16s, 32s, 64s, 128s, 256s, 512s, 1024s, 2048s, 4096s, 8192s, 16384s, -32768s, 0s, 0s, 0s, 0s, 0s, 0s, 0s, 0s, 0s, 0s, 0s, 0s, 0s, 0s ;
		Control_Flags_uncorr:flag_values = 2s, 4s, 8s, 16s, 32s, 64s, 128s, 256s, 512s, 1024s, 2048s, 4096s, 8192s, 16384s, -32768s, 0s, 0s, 0s, 0s, 0s, 0s, 0s, 0s, 0s, 0s, 0s, 0s, 0s, 0s ;
		string Control_Flags_uncorr:flag_meanings = "FG_CTRL_RANGE FG_CTRL_SIGMA FG_CTRL_CHI2 FG_CTRL_CHI2_P FG_CTRL_CONTAMINATED FG_CTRL_SUNGLINT FG_CTRL_MOONGLINT FG_CTRL_GAL_NOISE FG_CTRL_MIXED_SCENE FG_CTRL_REACH_MAXITER FG_CTRL_NUM_MEAS_MIN FG_CTRL_NUM_MEAS_LOW FG_CTRL_MANY_OUTLIERS FG_CTRL_MARQ FG_CTRL_ROUGHNESS FG_CTRL_FOAM FG_CTRL_ECMWF FG_CTRL_VALID FG_CTRL_NO_SURFACE FG_CTRL_RANGE_ACARD FG_CTRL_SIGMA_ACARD FG_CTRL_USED_FARATEC FG_CTRL_POOR_GEOPHYS FG_CTRL_POOR_RETRIEVAL FG_CTRL_SUSPECT_RFI FG_CTRL_RFI_PRONE_X FG_CTRL_RFI_PRONE_Y FG_CTRL_ADJUSTED_RA FG_CTRL_RETRIEV_FAIL" ;
		string Control_Flags_uncorr:_Unsigned = "true" ;
	ushort Dg_RFI_L1(n_grid_points) ;
		Dg_RFI_L1:_FillValue = 64537US ;
		string Dg_RFI_L1:_Unsigned = "true" ;
	ushort Dg_RFI_X(n_grid_points) ;
		Dg_RFI_X:_FillValue = 64537US ;
		string Dg_RFI_X:_Unsigned = "true" ;
	ushort Dg_RFI_Y(n_grid_points) ;
		Dg_RFI_Y:_FillValue = 64537US ;
		string Dg_RFI_Y:_Unsigned = "true" ;
	ushort Dg_RFI_probability(n_grid_points) ;
		string Dg_RFI_probability:units = "%" ;
		Dg_RFI_probability:_FillValue = 64537US ;
		string Dg_RFI_probability:_Unsigned = "true" ;
	ushort Dg_Suspect_ice(n_grid_points) ;
		Dg_Suspect_ice:_FillValue = 0US ;
		string Dg_Suspect_ice:_Unsigned = "true" ;
	ushort Dg_af_fov(n_grid_points) ;
		Dg_af_fov:_FillValue = 0US ;
		string Dg_af_fov:_Unsigned = "true" ;
	ushort Dg_border_fov(n_grid_points) ;
		Dg_border_fov:_FillValue = 0US ;
		string Dg_border_fov:_Unsigned = "true" ;
	ushort Dg_chi2_Acard(n_grid_points) ;
		Dg_chi2_Acard:_FillValue = 0US ;
		Dg_chi2_Acard:scale_factor = 0.00999999977648258 ;
		Dg_chi2_Acard:scale_offset = 0. ;
		string Dg_chi2_Acard:_Unsigned = "true" ;
	ushort Dg_chi2_P_Acard(n_grid_points) ;
		Dg_chi2_P_Acard:_FillValue = 0US ;
		Dg_chi2_P_Acard:scale_factor = 0.00100000004749745 ;
		Dg_chi2_P_Acard:scale_offset = 0. ;
		string Dg_chi2_P_Acard:_Unsigned = "true" ;
	ushort Dg_chi2_P_corr(n_grid_points) ;
		Dg_chi2_P_corr:_FillValue = 0US ;
		Dg_chi2_P_corr:scale_factor = 0.00100000004749745 ;
		Dg_chi2_P_corr:scale_offset = 0. ;
		string Dg_chi2_P_corr:_Unsigned = "true" ;
	ushort Dg_chi2_P_uncorr(n_grid_points) ;
		Dg_chi2_P_uncorr:_FillValue = 0US ;
		Dg_chi2_P_uncorr:scale_factor = 0.00100000004749745 ;
		Dg_chi2_P_uncorr:scale_offset = 0. ;
		string Dg_chi2_P_uncorr:_Unsigned = "true" ;
	ushort Dg_chi2_corr(n_grid_points) ;
		Dg_chi2_corr:_FillValue = 0US ;
		Dg_chi2_corr:scale_factor = 0.00999999977648258 ;
		Dg_chi2_corr:scale_offset = 0. ;
		string Dg_chi2_corr:_Unsigned = "true" ;
	ushort Dg_chi2_uncorr(n_grid_points) ;
		Dg_chi2_uncorr:_FillValue = 0US ;
		Dg_chi2_uncorr:scale_factor = 0.00999999977648258 ;
		Dg_chi2_uncorr:scale_offset = 0. ;
		string Dg_chi2_uncorr:_Unsigned = "true" ;
	ushort Dg_galactic_Noise_Error(n_grid_points) ;
		Dg_galactic_Noise_Error:_FillValue = 0US ;
		string Dg_galactic_Noise_Error:_Unsigned = "true" ;
	ushort Dg_moonglint(n_grid_points) ;
		Dg_moonglint:_FillValue = 0US ;
		string Dg_moonglint:_Unsigned = "true" ;
	ubyte Dg_num_iter_Acard(n_grid_points) ;
		Dg_num_iter_Acard:_FillValue = 0UB ;
		string Dg_num_iter_Acard:_Unsigned = "true" ;
	ubyte Dg_num_iter_corr(n_grid_points) ;
		Dg_num_iter_corr:_FillValue = 0UB ;
		string Dg_num_iter_corr:_Unsigned = "true" ;
	ubyte Dg_num_iter_uncorr(n_grid_points) ;
		Dg_num_iter_uncorr:_FillValue = 0UB ;
		string Dg_num_iter_uncorr:_Unsigned = "true" ;
	ushort Dg_num_meas_l1c(n_grid_points) ;
		Dg_num_meas_l1c:_FillValue = 0US ;
		string Dg_num_meas_l1c:_Unsigned = "true" ;
	ushort Dg_num_meas_valid(n_grid_points) ;
		Dg_num_meas_valid:_FillValue = 0US ;
		string Dg_num_meas_valid:_Unsigned = "true" ;
	ushort Dg_quality_SSS_anom(n_grid_points) ;
		Dg_quality_SSS_anom:_FillValue = 999US ;
		string Dg_quality_SSS_anom:_Unsigned = "true" ;
	ushort Dg_quality_SSS_corr(n_grid_points) ;
		Dg_quality_SSS_corr:_FillValue = 999US ;
		string Dg_quality_SSS_corr:_Unsigned = "true" ;
	ushort Dg_quality_SSS_uncorr(n_grid_points) ;
		Dg_quality_SSS_uncorr:_FillValue = 999US ;
		string Dg_quality_SSS_uncorr:_Unsigned = "true" ;
	ushort Dg_sky(n_grid_points) ;
		Dg_sky:_FillValue = 64537US ;
		string Dg_sky:_Unsigned = "true" ;
	ushort Dg_sun_glint_L2(n_grid_points) ;
		Dg_sun_glint_L2:_FillValue = 0US ;
		string Dg_sun_glint_L2:_Unsigned = "true" ;
	ushort Dg_sun_glint_area(n_grid_points) ;
		Dg_sun_glint_area:_FillValue = 0US ;
		string Dg_sun_glint_area:_Unsigned = "true" ;
	ushort Dg_sun_glint_fov(n_grid_points) ;
		Dg_sun_glint_fov:_FillValue = 0US ;
		string Dg_sun_glint_fov:_Unsigned = "true" ;
	ushort Dg_sun_tails(n_grid_points) ;
		Dg_sun_tails:_FillValue = 0US ;
		string Dg_sun_tails:_Unsigned = "true" ;
	float Equiv_ftprt_diam(n_grid_points) ;
		string Equiv_ftprt_diam:units = "km" ;
		Equiv_ftprt_diam:_FillValue = -999.f ;
	uint Grid_Point_ID(n_grid_points) ;
		Grid_Point_ID:_FillValue = 0U ;
		string Grid_Point_ID:_Unsigned = "true" ;
	float Latitude(n_grid_points) ;
		string Latitude:units = "deg" ;
		Latitude:_FillValue = -999.f ;
	float Longitude(n_grid_points) ;
		string Longitude:units = "deg" ;
		Longitude:_FillValue = -999.f ;
	float Mean_acq_time(n_grid_points) ;
		string Mean_acq_time:units = "dd" ;
		Mean_acq_time:_FillValue = -999.f ;
	float SSS_anom(n_grid_points) ;
		string SSS_anom:units = "psu" ;
		SSS_anom:_FillValue = -999.f ;
	ushort SSS_climatology(n_grid_points) ;
		SSS_climatology:_FillValue = 0US ;
		SSS_climatology:scale_factor = 0.00999999977648258 ;
		SSS_climatology:scale_offset = 0. ;
		string SSS_climatology:_Unsigned = "true" ;
	float SSS_corr(n_grid_points) ;
		string SSS_corr:units = "psu" ;
		SSS_corr:_FillValue = -999.f ;
	float SSS_uncorr(n_grid_points) ;
		string SSS_uncorr:units = "psu" ;
		SSS_uncorr:_FillValue = -999.f ;
	float SST(n_grid_points) ;
		string SST:units = "°C" ;
		SST:_FillValue = -999.f ;
	uint Science_Flags_Acard(n_grid_points) ;
		Science_Flags_Acard:_FillValue = 0U ;
		Science_Flags_Acard:flag_masks = 1s, 2s, 4s, 8s, 16s, 32s, 64s, 128s, 256s, 512s, 1024s, 2048s, 4096s, 8192s, 16384s, -32768s, 0s, 0s, 0s, 0s, 0s, 0s, 0s ;
		Science_Flags_Acard:flag_values = 1s, 2s, 4s, 8s, 16s, 32s, 64s, 128s, 256s, 512s, 1024s, 2048s, 4096s, 8192s, 16384s, -32768s, 0s, 0s, 0s, 0s, 0s, 0s, 0s ;
		string Science_Flags_Acard:flag_meanings = "FG_SC_LAND_SEA_COAST1 FG_SC_LAND_SEA_COAST2 FG_SC_TEC_GRADIENT FG_SC_IN_CLIM_ICE FG_SC_ICE FG_SC_SUSPECT_ICE FG_SC_RAIN FG_SC_HIGH_WIND FG_SC_LOW_WIND FG_SC_HIGHT_SST FG_SC_LOW_SST FG_SC_HIGH_SSS FG_SC_LOW_SSS FG_SC_SEA_STATE_1 FG_SC_SEA_STATE_2 FG_SC_SEA_STATE_3 FG_SC_SEA_STATE_4 FG_SC_SEA_STATE_5 FG_SC_SEA_STATE_6 FG_SC_SST_FRONT FG_SC_SSS_FRONT FG_SC_ICE_ACARD FG_SC_ECMWF_LAND" ;
		string Science_Flags_Acard:_Unsigned = "true" ;
	uint Science_Flags_anom(n_grid_points) ;
		Science_Flags_anom:_FillValue = 0U ;
		Science_Flags_anom:flag_masks = 1s, 2s, 4s, 8s, 16s, 32s, 64s, 128s, 256s, 512s, 1024s, 2048s, 4096s, 8192s, 16384s, -32768s, 0s, 0s, 0s, 0s, 0s, 0s, 0s ;
		Science_Flags_anom:flag_values = 1s, 2s, 4s, 8s, 16s, 32s, 64s, 128s, 256s, 512s, 1024s, 2048s, 4096s, 8192s, 16384s, -32768s, 0s, 0s, 0s, 0s, 0s, 0s, 0s ;
		string Science_Flags_anom:flag_meanings = "FG_SC_LAND_SEA_COAST1 FG_SC_LAND_SEA_COAST2 FG_SC_TEC_GRADIENT FG_SC_IN_CLIM_ICE FG_SC_ICE FG_SC_SUSPECT_ICE FG_SC_RAIN FG_SC_HIGH_WIND FG_SC_LOW_WIND FG_SC_HIGHT_SST FG_SC_LOW_SST FG_SC_HIGH_SSS FG_SC_LOW_SSS FG_SC_SEA_STATE_1 FG_SC_SEA_STATE_2 FG_SC_SEA_STATE_3 FG_SC_SEA_STATE_4 FG_SC_SEA_STATE_5 FG_SC_SEA_STATE_6 FG_SC_SST_FRONT FG_SC_SSS_FRONT FG_SC_ICE_ACARD FG_SC_ECMWF_LAND" ;
		string Science_Flags_anom:_Unsigned = "true" ;
	uint Science_Flags_corr(n_grid_points) ;
		Science_Flags_corr:_FillValue = 0U ;
		Science_Flags_corr:flag_masks = 1s, 2s, 4s, 8s, 16s, 32s, 64s, 128s, 256s, 512s, 1024s, 2048s, 4096s, 8192s, 16384s, -32768s, 0s, 0s, 0s, 0s, 0s, 0s, 0s ;
		Science_Flags_corr:flag_values = 1s, 2s, 4s, 8s, 16s, 32s, 64s, 128s, 256s, 512s, 1024s, 2048s, 4096s, 8192s, 16384s, -32768s, 0s, 0s, 0s, 0s, 0s, 0s, 0s ;
		string Science_Flags_corr:flag_meanings = "FG_SC_LAND_SEA_COAST1 FG_SC_LAND_SEA_COAST2 FG_SC_TEC_GRADIENT FG_SC_IN_CLIM_ICE FG_SC_ICE FG_SC_SUSPECT_ICE FG_SC_RAIN FG_SC_HIGH_WIND FG_SC_LOW_WIND FG_SC_HIGHT_SST FG_SC_LOW_SST FG_SC_HIGH_SSS FG_SC_LOW_SSS FG_SC_SEA_STATE_1 FG_SC_SEA_STATE_2 FG_SC_SEA_STATE_3 FG_SC_SEA_STATE_4 FG_SC_SEA_STATE_5 FG_SC_SEA_STATE_6 FG_SC_SST_FRONT FG_SC_SSS_FRONT FG_SC_ICE_ACARD FG_SC_ECMWF_LAND" ;
		string Science_Flags_corr:_Unsigned = "true" ;
	uint Science_Flags_uncorr(n_grid_points) ;
		Science_Flags_uncorr:_FillValue = 0U ;
		Science_Flags_uncorr:flag_masks = 1s, 2s, 4s, 8s, 16s, 32s, 64s, 128s, 256s, 512s, 1024s, 2048s, 4096s, 8192s, 16384s, -32768s, 0s, 0s, 0s, 0s, 0s, 0s, 0s ;
		Science_Flags_uncorr:flag_values = 1s, 2s, 4s, 8s, 16s, 32s, 64s, 128s, 256s, 512s, 1024s, 2048s, 4096s, 8192s, 16384s, -32768s, 0s, 0s, 0s, 0s, 0s, 0s, 0s ;
		string Science_Flags_uncorr:flag_meanings = "FG_SC_LAND_SEA_COAST1 FG_SC_LAND_SEA_COAST2 FG_SC_TEC_GRADIENT FG_SC_IN_CLIM_ICE FG_SC_ICE FG_SC_SUSPECT_ICE FG_SC_RAIN FG_SC_HIGH_WIND FG_SC_LOW_WIND FG_SC_HIGHT_SST FG_SC_LOW_SST FG_SC_HIGH_SSS FG_SC_LOW_SSS FG_SC_SEA_STATE_1 FG_SC_SEA_STATE_2 FG_SC_SEA_STATE_3 FG_SC_SEA_STATE_4 FG_SC_SEA_STATE_5 FG_SC_SEA_STATE_6 FG_SC_SST_FRONT FG_SC_SSS_FRONT FG_SC_ICE_ACARD FG_SC_ECMWF_LAND" ;
		string Science_Flags_uncorr:_Unsigned = "true" ;
	float Sigma_Acard(n_grid_points) ;
		Sigma_Acard:_FillValue = -999.f ;
	float Sigma_SSS_anom(n_grid_points) ;
		string Sigma_SSS_anom:units = "psu" ;
		Sigma_SSS_anom:_FillValue = -999.f ;
	float Sigma_SSS_corr(n_grid_points) ;
		string Sigma_SSS_corr:units = "psu" ;
		Sigma_SSS_corr:_FillValue = -999.f ;
	float Sigma_SSS_uncorr(n_grid_points) ;
		string Sigma_SSS_uncorr:units = "psu" ;
		Sigma_SSS_uncorr:_FillValue = -999.f ;
	float Sigma_Tb_42_5H(n_grid_points) ;
		string Sigma_Tb_42_5H:units = "K" ;
		Sigma_Tb_42_5H:_FillValue = -999.f ;
	float Sigma_Tb_42_5V(n_grid_points) ;
		string Sigma_Tb_42_5V:units = "K" ;
		Sigma_Tb_42_5V:_FillValue = -999.f ;
	float Sigma_Tb_42_5X(n_grid_points) ;
		string Sigma_Tb_42_5X:units = "K" ;
		Sigma_Tb_42_5X:_FillValue = -999.f ;
	float Sigma_Tb_42_5Y(n_grid_points) ;
		string Sigma_Tb_42_5Y:units = "K" ;
		Sigma_Tb_42_5Y:_FillValue = -999.f ;
	ushort Sigma_WS_corr(n_grid_points) ;
		Sigma_WS_corr:_FillValue = 0US ;
		Sigma_WS_corr:scale_factor = 0.00100000004749745 ;
		Sigma_WS_corr:scale_offset = 0. ;
		string Sigma_WS_corr:_Unsigned = "true" ;
	float Tb_42_5H(n_grid_points) ;
		string Tb_42_5H:units = "K" ;
		Tb_42_5H:_FillValue = -999.f ;
	float Tb_42_5V(n_grid_points) ;
		string Tb_42_5V:units = "K" ;
		Tb_42_5V:_FillValue = -999.f ;
	float Tb_42_5X(n_grid_points) ;
		string Tb_42_5X:units = "K" ;
		Tb_42_5X:_FillValue = -999.f ;
	float Tb_42_5Y(n_grid_points) ;
		string Tb_42_5Y:units = "K" ;
		Tb_42_5Y:_FillValue = -999.f ;
	float WS(n_grid_points) ;
		string WS:units = "m s-1" ;
		WS:_FillValue = -999.f ;
	ushort WS_corr(n_grid_points) ;
		WS_corr:_FillValue = 0US ;
		WS_corr:scale_factor = 0.00100000004749745 ;
		WS_corr:scale_offset = 0. ;
		string WS_corr:_Unsigned = "true" ;
	float X_swath(n_grid_points) ;
		string X_swath:units = "m" ;
		X_swath:_FillValue = -999.f ;

// global attributes:
		string :creation_date = "UTC=2021-07-01T05:16:26" ;
		string :total_number_of_grid_points = "92713" ;
		string :FH\:File_Name = "SM_OPER_MIR_OSUDP2_20210630T215911_20210630T225230_700_001_1" ;
		string :FH\:File_Description = "L2 Ocean Salinity Output User Data Product." ;
		string :FH\:Notes = "The UDP (User Data Product) is designed for oceanographics and high level centers, it includes geophysical parameters, a theoretical estimate of their accuracy, flags and descriptors of the product quality." ;
		string :FH\:Mission = "SMOS" ;
		string :FH\:File_Class = "OPER" ;
		string :FH\:File_Type = "MIR_OSUDP2" ;
		string :FH\:File_Version = "0001" ;
		string :FH\:Validity_Period\:Validity_Start = "UTC=2021-06-30T21:59:11" ;
		string :FH\:Validity_Period\:Validity_Stop = "UTC=2021-06-30T22:52:30" ;
		string :FH\:Source\:System = "DPGS" ;
		string :FH\:Source\:Creator = "L2OP" ;
		string :FH\:Source\:Creator_Version = "700" ;
		string :FH\:Source\:Creation_Date = "UTC=2021-07-01T05:09:30" ;
		string :VH\:SPH\:QI\:Total_Selected_L1c_Grid_Points = "60219" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:Retrieval_Scheme = "1" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:Land_Rejected = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:Too_Close_To_Land_Rejected = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:Ice_Rejected = "10855" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:Missing_ECMWF_Rejected = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:Too_Few_Measurements_Rejected = "18084" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:Good_Quality_Grid_Points = "29636" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:Poor_Quality_Grid_Points = "4896" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:SQ\:Grid_Point_Type = "Sea" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:SQ\:SSS_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:SQ\:SST_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:SQ\:WS_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:SQ\:Good_Quality = "23293" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:SQ\:Good_Quality_Retrieved = "17816" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:SQ\:Good_Quality_Retrieved_Average_Sigma = "1.959542" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:SQ\:Good_Quality_Failed_Outside_Valid_Range = "81" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:SQ\:Good_Quality_Failed_Sigma_Too_High = "478" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:SQ\:Good_Quality_Failed_Poor_Fit = "5037" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:SQ\:Good_Quality_Failed_Marquardt = "4" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:SQ\:Good_Quality_Failed_Maxiter = "110" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:SQ\:Good_Quality_Failed_OOLUT = "555" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:SQ\:Poor_Quality = "2426" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:SQ\:Poor_Quality_Retrieved = "1661" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:SQ\:Poor_Quality_Retrieved_Average_Sigma = "2.933723" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:NCQ\:Grid_Point_Type = "Near_Coast" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:NCQ\:SSS_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:NCQ\:SST_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:NCQ\:WS_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:NCQ\:Good_Quality = "6343" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:NCQ\:Good_Quality_Retrieved = "3803" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:NCQ\:Good_Quality_Retrieved_Average_Sigma = "1.253443" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:NCQ\:Good_Quality_Failed_Outside_Valid_Range = "276" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:NCQ\:Good_Quality_Failed_Sigma_Too_High = "522" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:NCQ\:Good_Quality_Failed_Poor_Fit = "2247" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:NCQ\:Good_Quality_Failed_Marquardt = "152" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:NCQ\:Good_Quality_Failed_Maxiter = "411" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:NCQ\:Good_Quality_Failed_OOLUT = "773" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:NCQ\:Poor_Quality = "2470" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:NCQ\:Poor_Quality_Retrieved = "1367" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:NCQ\:Poor_Quality_Retrieved_Average_Sigma = "1.480500" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_0\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_0\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_0\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_0\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_0\:Good_Quality = "559" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_0\:Good_Quality_Retrieved = "131" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_0\:Good_Quality_Retrieved_Average_Sigma = "1.985529" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_0\:Good_Quality_Failed_Outside_Valid_Range = "183" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_0\:Good_Quality_Failed_Sigma_Too_High = "261" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_0\:Good_Quality_Failed_Poor_Fit = "325" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_0\:Good_Quality_Failed_Marquardt = "112" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_0\:Good_Quality_Failed_Maxiter = "130" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_0\:Good_Quality_Failed_OOLUT = "326" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_0\:Poor_Quality = "106" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_0\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_0\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_1\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_1\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_1\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_1\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_1\:Good_Quality = "486" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_1\:Good_Quality_Retrieved = "229" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_1\:Good_Quality_Retrieved_Average_Sigma = "2.167454" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_1\:Good_Quality_Failed_Outside_Valid_Range = "60" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_1\:Good_Quality_Failed_Sigma_Too_High = "82" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_1\:Good_Quality_Failed_Poor_Fit = "244" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_1\:Good_Quality_Failed_Marquardt = "30" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_1\:Good_Quality_Failed_Maxiter = "45" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_1\:Good_Quality_Failed_OOLUT = "135" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_1\:Poor_Quality = "233" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_1\:Poor_Quality_Retrieved = "13" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_1\:Poor_Quality_Retrieved_Average_Sigma = "4.597799" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_2\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_2\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_2\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_2\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_2\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_2\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_2\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_2\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_2\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_2\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_2\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_2\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_2\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_2\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_2\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_2\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_3\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_3\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_3\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_3\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_3\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_3\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_3\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_3\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_3\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_3\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_3\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_3\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_3\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_3\:Poor_Quality = "3" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_3\:Poor_Quality_Retrieved = "1" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_3\:Poor_Quality_Retrieved_Average_Sigma = "2.726585" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_4\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_4\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_4\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_4\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_4\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_4\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_4\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_4\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_4\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_4\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_4\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_4\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_4\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_4\:Poor_Quality = "233" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_4\:Poor_Quality_Retrieved = "182" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_4\:Poor_Quality_Retrieved_Average_Sigma = "3.945308" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_5\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_5\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_5\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_5\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_5\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_5\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_5\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_5\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_5\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_5\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_5\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_5\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_5\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_5\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_5\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_5\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_6\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_6\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_6\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_6\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_6\:Good_Quality = "16" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_6\:Good_Quality_Retrieved = "14" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_6\:Good_Quality_Retrieved_Average_Sigma = "1.307737" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_6\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_6\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_6\:Good_Quality_Failed_Poor_Fit = "2" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_6\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_6\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_6\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_6\:Poor_Quality = "22" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_6\:Poor_Quality_Retrieved = "19" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_6\:Poor_Quality_Retrieved_Average_Sigma = "1.902701" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_7\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_7\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_7\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_7\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_7\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_7\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_7\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_7\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_7\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_7\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_7\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_7\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_7\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_7\:Poor_Quality = "113" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_7\:Poor_Quality_Retrieved = "58" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_7\:Poor_Quality_Retrieved_Average_Sigma = "1.925949" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_8\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_8\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_8\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_8\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_8\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_8\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_8\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_8\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_8\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_8\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_8\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_8\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_8\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_8\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_8\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_8\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_9\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_9\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_9\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_9\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_9\:Good_Quality = "1485" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_9\:Good_Quality_Retrieved = "825" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_9\:Good_Quality_Retrieved_Average_Sigma = "2.191673" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_9\:Good_Quality_Failed_Outside_Valid_Range = "1" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_9\:Good_Quality_Failed_Sigma_Too_High = "54" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_9\:Good_Quality_Failed_Poor_Fit = "544" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_9\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_9\:Good_Quality_Failed_Maxiter = "247" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_9\:Good_Quality_Failed_OOLUT = "190" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_9\:Poor_Quality = "11" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_9\:Poor_Quality_Retrieved = "1" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_9\:Poor_Quality_Retrieved_Average_Sigma = "4.534814" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_10\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_10\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_10\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_10\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_10\:Good_Quality = "6940" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_10\:Good_Quality_Retrieved = "4685" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_10\:Good_Quality_Retrieved_Average_Sigma = "2.611991" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_10\:Good_Quality_Failed_Outside_Valid_Range = "102" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_10\:Good_Quality_Failed_Sigma_Too_High = "600" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_10\:Good_Quality_Failed_Poor_Fit = "1779" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_10\:Good_Quality_Failed_Marquardt = "14" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_10\:Good_Quality_Failed_Maxiter = "72" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_10\:Good_Quality_Failed_OOLUT = "603" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_10\:Poor_Quality = "508" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_10\:Poor_Quality_Retrieved = "218" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_10\:Poor_Quality_Retrieved_Average_Sigma = "4.334874" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_11\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_11\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_11\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_11\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_11\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_11\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_11\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_11\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_11\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_11\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_11\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_11\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_11\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_11\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_11\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_11\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_12\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_12\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_12\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_12\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_12\:Good_Quality = "232" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_12\:Good_Quality_Retrieved = "156" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_12\:Good_Quality_Retrieved_Average_Sigma = "1.521774" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_12\:Good_Quality_Failed_Outside_Valid_Range = "1" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_12\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_12\:Good_Quality_Failed_Poor_Fit = "70" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_12\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_12\:Good_Quality_Failed_Maxiter = "7" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_12\:Good_Quality_Failed_OOLUT = "17" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_12\:Poor_Quality = "55" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_12\:Poor_Quality_Retrieved = "42" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_12\:Poor_Quality_Retrieved_Average_Sigma = "2.482193" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_13\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_13\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_13\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_13\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_13\:Good_Quality = "11990" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_13\:Good_Quality_Retrieved = "9532" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_13\:Good_Quality_Retrieved_Average_Sigma = "2.064730" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_13\:Good_Quality_Failed_Outside_Valid_Range = "10" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_13\:Good_Quality_Failed_Sigma_Too_High = "3" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_13\:Good_Quality_Failed_Poor_Fit = "2454" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_13\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_13\:Good_Quality_Failed_Maxiter = "1" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_13\:Good_Quality_Failed_OOLUT = "42" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_13\:Poor_Quality = "997" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_13\:Poor_Quality_Retrieved = "857" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_13\:Poor_Quality_Retrieved_Average_Sigma = "3.092174" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_14\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_14\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_14\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_14\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_14\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_14\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_14\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_14\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_14\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_14\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_14\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_14\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_14\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_14\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_14\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_14\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_15\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_15\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_15\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_15\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_15\:Good_Quality = "830" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_15\:Good_Quality_Retrieved = "677" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_15\:Good_Quality_Retrieved_Average_Sigma = "1.047869" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_15\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_15\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_15\:Good_Quality_Failed_Poor_Fit = "153" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_15\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_15\:Good_Quality_Failed_Maxiter = "1" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_15\:Good_Quality_Failed_OOLUT = "4" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_15\:Poor_Quality = "1379" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_15\:Poor_Quality_Retrieved = "1092" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_15\:Poor_Quality_Retrieved_Average_Sigma = "1.087475" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_16\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_16\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_16\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_16\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_16\:Good_Quality = "7097" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_16\:Good_Quality_Retrieved = "5369" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_16\:Good_Quality_Retrieved_Average_Sigma = "0.787403" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_16\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_16\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_16\:Good_Quality_Failed_Poor_Fit = "1713" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_16\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_16\:Good_Quality_Failed_Maxiter = "18" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_16\:Good_Quality_Failed_OOLUT = "11" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_16\:Poor_Quality = "1043" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_16\:Poor_Quality_Retrieved = "450" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_16\:Poor_Quality_Retrieved_Average_Sigma = "1.581808" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_17\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_17\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_17\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_17\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_17\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_17\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_17\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_17\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_17\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_17\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_17\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_17\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_17\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_17\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_17\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_17\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_18\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_18\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_18\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_18\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_18\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_18\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_18\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_18\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_18\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_18\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_18\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_18\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_18\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_18\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_18\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_18\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_19\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_19\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_19\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_19\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_19\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_19\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_19\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_19\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_19\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_19\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_19\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_19\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_19\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_19\:Poor_Quality = "141" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_19\:Poor_Quality_Retrieved = "51" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_19\:Poor_Quality_Retrieved_Average_Sigma = "4.372903" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_20\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_20\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_20\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_20\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_20\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_20\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_20\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_20\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_20\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_20\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_20\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_20\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_20\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_20\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_20\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_20\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_21\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_21\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_21\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_21\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_21\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_21\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_21\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_21\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_21\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_21\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_21\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_21\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_21\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_21\:Poor_Quality = "8" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_21\:Poor_Quality_Retrieved = "5" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_21\:Poor_Quality_Retrieved_Average_Sigma = "2.769263" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_22\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_22\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_22\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_22\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_22\:Good_Quality = "1" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_22\:Good_Quality_Retrieved = "1" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_22\:Good_Quality_Retrieved_Average_Sigma = "2.597888" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_22\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_22\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_22\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_22\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_22\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_22\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_22\:Poor_Quality = "42" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_22\:Poor_Quality_Retrieved = "37" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_22\:Poor_Quality_Retrieved_Average_Sigma = "3.355307" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_23\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_23\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_23\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_23\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_23\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_23\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_23\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_23\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_23\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_23\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_23\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_23\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_23\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_23\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_23\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_23\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_24\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_24\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_24\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_24\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_24\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_24\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_24\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_24\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_24\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_24\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_24\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_24\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_24\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_24\:Poor_Quality = "2" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_24\:Poor_Quality_Retrieved = "2" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_24\:Poor_Quality_Retrieved_Average_Sigma = "2.113266" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_25\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_25\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_25\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_25\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_25\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_25\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_25\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_25\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_25\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_25\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_25\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_25\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_25\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_25\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_25\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_25\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_26\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_26\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_26\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_26\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_26\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_26\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_26\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_26\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_26\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_26\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_26\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_26\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_26\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_26\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_26\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_26\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:SIQ\:Grid_Point_Type = "Sea_Ice" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:SIQ\:SSS_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:SIQ\:SST_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:SIQ\:WS_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:SIQ\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:SIQ\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:SIQ\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:SIQ\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:SIQ\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:SIQ\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:SIQ\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:SIQ\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:SIQ\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:SIQ\:Poor_Quality = "64" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:SIQ\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:SIQ\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:Retrieval_Scheme = "2" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:Land_Rejected = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:Too_Close_To_Land_Rejected = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:Ice_Rejected = "10855" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:Missing_ECMWF_Rejected = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:Too_Few_Measurements_Rejected = "18084" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:Good_Quality_Grid_Points = "29636" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:Poor_Quality_Grid_Points = "4896" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:SQ\:Grid_Point_Type = "Sea" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:SQ\:SSS_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:SQ\:SST_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:SQ\:WS_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:SQ\:Good_Quality = "23293" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:SQ\:Good_Quality_Retrieved = "16753" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:SQ\:Good_Quality_Retrieved_Average_Sigma = "2.016282" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:SQ\:Good_Quality_Failed_Outside_Valid_Range = "78" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:SQ\:Good_Quality_Failed_Sigma_Too_High = "479" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:SQ\:Good_Quality_Failed_Poor_Fit = "5999" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:SQ\:Good_Quality_Failed_Marquardt = "4" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:SQ\:Good_Quality_Failed_Maxiter = "273" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:SQ\:Good_Quality_Failed_OOLUT = "555" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:SQ\:Poor_Quality = "2426" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:SQ\:Poor_Quality_Retrieved = "1638" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:SQ\:Poor_Quality_Retrieved_Average_Sigma = "2.984403" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:NCQ\:Grid_Point_Type = "Near_Coast" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:NCQ\:SSS_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:NCQ\:SST_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:NCQ\:WS_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:NCQ\:Good_Quality = "6343" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:NCQ\:Good_Quality_Retrieved = "2879" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:NCQ\:Good_Quality_Retrieved_Average_Sigma = "1.380678" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:NCQ\:Good_Quality_Failed_Outside_Valid_Range = "281" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:NCQ\:Good_Quality_Failed_Sigma_Too_High = "532" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:NCQ\:Good_Quality_Failed_Poor_Fit = "3163" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:NCQ\:Good_Quality_Failed_Marquardt = "167" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:NCQ\:Good_Quality_Failed_Maxiter = "402" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:NCQ\:Good_Quality_Failed_OOLUT = "818" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:NCQ\:Poor_Quality = "2470" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:NCQ\:Poor_Quality_Retrieved = "1286" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:NCQ\:Poor_Quality_Retrieved_Average_Sigma = "1.503417" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_0\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_0\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_0\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_0\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_0\:Good_Quality = "559" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_0\:Good_Quality_Retrieved = "130" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_0\:Good_Quality_Retrieved_Average_Sigma = "1.956271" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_0\:Good_Quality_Failed_Outside_Valid_Range = "189" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_0\:Good_Quality_Failed_Sigma_Too_High = "265" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_0\:Good_Quality_Failed_Poor_Fit = "323" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_0\:Good_Quality_Failed_Marquardt = "121" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_0\:Good_Quality_Failed_Maxiter = "121" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_0\:Good_Quality_Failed_OOLUT = "326" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_0\:Poor_Quality = "106" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_0\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_0\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_1\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_1\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_1\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_1\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_1\:Good_Quality = "486" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_1\:Good_Quality_Retrieved = "228" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_1\:Good_Quality_Retrieved_Average_Sigma = "2.158294" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_1\:Good_Quality_Failed_Outside_Valid_Range = "59" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_1\:Good_Quality_Failed_Sigma_Too_High = "85" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_1\:Good_Quality_Failed_Poor_Fit = "245" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_1\:Good_Quality_Failed_Marquardt = "36" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_1\:Good_Quality_Failed_Maxiter = "40" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_1\:Good_Quality_Failed_OOLUT = "136" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_1\:Poor_Quality = "233" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_1\:Poor_Quality_Retrieved = "13" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_1\:Poor_Quality_Retrieved_Average_Sigma = "4.621669" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_2\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_2\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_2\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_2\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_2\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_2\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_2\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_2\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_2\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_2\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_2\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_2\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_2\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_2\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_2\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_2\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_3\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_3\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_3\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_3\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_3\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_3\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_3\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_3\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_3\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_3\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_3\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_3\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_3\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_3\:Poor_Quality = "3" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_3\:Poor_Quality_Retrieved = "1" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_3\:Poor_Quality_Retrieved_Average_Sigma = "2.825164" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_4\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_4\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_4\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_4\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_4\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_4\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_4\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_4\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_4\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_4\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_4\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_4\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_4\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_4\:Poor_Quality = "233" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_4\:Poor_Quality_Retrieved = "182" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_4\:Poor_Quality_Retrieved_Average_Sigma = "4.031709" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_5\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_5\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_5\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_5\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_5\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_5\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_5\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_5\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_5\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_5\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_5\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_5\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_5\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_5\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_5\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_5\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_6\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_6\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_6\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_6\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_6\:Good_Quality = "16" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_6\:Good_Quality_Retrieved = "14" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_6\:Good_Quality_Retrieved_Average_Sigma = "1.316742" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_6\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_6\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_6\:Good_Quality_Failed_Poor_Fit = "2" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_6\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_6\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_6\:Good_Quality_Failed_OOLUT = "1" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_6\:Poor_Quality = "22" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_6\:Poor_Quality_Retrieved = "16" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_6\:Poor_Quality_Retrieved_Average_Sigma = "1.820999" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_7\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_7\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_7\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_7\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_7\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_7\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_7\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_7\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_7\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_7\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_7\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_7\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_7\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_7\:Poor_Quality = "113" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_7\:Poor_Quality_Retrieved = "48" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_7\:Poor_Quality_Retrieved_Average_Sigma = "1.882463" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_8\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_8\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_8\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_8\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_8\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_8\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_8\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_8\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_8\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_8\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_8\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_8\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_8\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_8\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_8\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_8\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_9\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_9\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_9\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_9\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_9\:Good_Quality = "1485" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_9\:Good_Quality_Retrieved = "821" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_9\:Good_Quality_Retrieved_Average_Sigma = "2.183326" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_9\:Good_Quality_Failed_Outside_Valid_Range = "2" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_9\:Good_Quality_Failed_Sigma_Too_High = "57" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_9\:Good_Quality_Failed_Poor_Fit = "544" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_9\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_9\:Good_Quality_Failed_Maxiter = "247" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_9\:Good_Quality_Failed_OOLUT = "194" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_9\:Poor_Quality = "11" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_9\:Poor_Quality_Retrieved = "1" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_9\:Poor_Quality_Retrieved_Average_Sigma = "4.586421" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_10\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_10\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_10\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_10\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_10\:Good_Quality = "6940" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_10\:Good_Quality_Retrieved = "4685" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_10\:Good_Quality_Retrieved_Average_Sigma = "2.610784" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_10\:Good_Quality_Failed_Outside_Valid_Range = "102" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_10\:Good_Quality_Failed_Sigma_Too_High = "601" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_10\:Good_Quality_Failed_Poor_Fit = "1779" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_10\:Good_Quality_Failed_Marquardt = "14" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_10\:Good_Quality_Failed_Maxiter = "71" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_10\:Good_Quality_Failed_OOLUT = "604" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_10\:Poor_Quality = "508" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_10\:Poor_Quality_Retrieved = "216" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_10\:Poor_Quality_Retrieved_Average_Sigma = "4.321773" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_11\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_11\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_11\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_11\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_11\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_11\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_11\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_11\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_11\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_11\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_11\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_11\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_11\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_11\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_11\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_11\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_12\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_12\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_12\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_12\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_12\:Good_Quality = "232" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_12\:Good_Quality_Retrieved = "154" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_12\:Good_Quality_Retrieved_Average_Sigma = "1.546095" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_12\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_12\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_12\:Good_Quality_Failed_Poor_Fit = "73" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_12\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_12\:Good_Quality_Failed_Maxiter = "5" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_12\:Good_Quality_Failed_OOLUT = "17" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_12\:Poor_Quality = "55" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_12\:Poor_Quality_Retrieved = "44" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_12\:Poor_Quality_Retrieved_Average_Sigma = "2.515923" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_13\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_13\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_13\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_13\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_13\:Good_Quality = "11990" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_13\:Good_Quality_Retrieved = "9022" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_13\:Good_Quality_Retrieved_Average_Sigma = "2.096603" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_13\:Good_Quality_Failed_Outside_Valid_Range = "7" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_13\:Good_Quality_Failed_Sigma_Too_High = "3" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_13\:Good_Quality_Failed_Poor_Fit = "2966" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_13\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_13\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_13\:Good_Quality_Failed_OOLUT = "58" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_13\:Poor_Quality = "997" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_13\:Poor_Quality_Retrieved = "849" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_13\:Poor_Quality_Retrieved_Average_Sigma = "3.150212" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_14\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_14\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_14\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_14\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_14\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_14\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_14\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_14\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_14\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_14\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_14\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_14\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_14\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_14\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_14\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_14\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_15\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_15\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_15\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_15\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_15\:Good_Quality = "830" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_15\:Good_Quality_Retrieved = "539" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_15\:Good_Quality_Retrieved_Average_Sigma = "1.062494" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_15\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_15\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_15\:Good_Quality_Failed_Poor_Fit = "288" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_15\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_15\:Good_Quality_Failed_Maxiter = "3" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_15\:Good_Quality_Failed_OOLUT = "13" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_15\:Poor_Quality = "1379" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_15\:Poor_Quality_Retrieved = "1021" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_15\:Poor_Quality_Retrieved_Average_Sigma = "1.095964" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_16\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_16\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_16\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_16\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_16\:Good_Quality = "7097" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_16\:Good_Quality_Retrieved = "4038" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_16\:Good_Quality_Retrieved_Average_Sigma = "0.801339" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_16\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_16\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_16\:Good_Quality_Failed_Poor_Fit = "2942" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_16\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_16\:Good_Quality_Failed_Maxiter = "188" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_16\:Good_Quality_Failed_OOLUT = "24" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_16\:Poor_Quality = "1043" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_16\:Poor_Quality_Retrieved = "438" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_16\:Poor_Quality_Retrieved_Average_Sigma = "1.589996" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_17\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_17\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_17\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_17\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_17\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_17\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_17\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_17\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_17\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_17\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_17\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_17\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_17\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_17\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_17\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_17\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_18\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_18\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_18\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_18\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_18\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_18\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_18\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_18\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_18\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_18\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_18\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_18\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_18\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_18\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_18\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_18\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_19\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_19\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_19\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_19\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_19\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_19\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_19\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_19\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_19\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_19\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_19\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_19\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_19\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_19\:Poor_Quality = "141" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_19\:Poor_Quality_Retrieved = "52" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_19\:Poor_Quality_Retrieved_Average_Sigma = "4.370056" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_20\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_20\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_20\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_20\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_20\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_20\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_20\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_20\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_20\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_20\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_20\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_20\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_20\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_20\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_20\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_20\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_21\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_21\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_21\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_21\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_21\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_21\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_21\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_21\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_21\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_21\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_21\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_21\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_21\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_21\:Poor_Quality = "8" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_21\:Poor_Quality_Retrieved = "5" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_21\:Poor_Quality_Retrieved_Average_Sigma = "2.781770" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_22\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_22\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_22\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_22\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_22\:Good_Quality = "1" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_22\:Good_Quality_Retrieved = "1" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_22\:Good_Quality_Retrieved_Average_Sigma = "2.728715" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_22\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_22\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_22\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_22\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_22\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_22\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_22\:Poor_Quality = "42" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_22\:Poor_Quality_Retrieved = "36" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_22\:Poor_Quality_Retrieved_Average_Sigma = "3.373684" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_23\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_23\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_23\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_23\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_23\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_23\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_23\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_23\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_23\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_23\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_23\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_23\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_23\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_23\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_23\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_23\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_24\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_24\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_24\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_24\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_24\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_24\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_24\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_24\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_24\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_24\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_24\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_24\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_24\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_24\:Poor_Quality = "2" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_24\:Poor_Quality_Retrieved = "2" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_24\:Poor_Quality_Retrieved_Average_Sigma = "2.176347" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_25\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_25\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_25\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_25\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_25\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_25\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_25\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_25\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_25\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_25\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_25\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_25\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_25\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_25\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_25\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_25\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_26\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_26\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_26\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_26\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_26\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_26\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_26\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_26\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_26\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_26\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_26\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_26\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_26\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_26\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_26\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_26\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:SIQ\:Grid_Point_Type = "Sea_Ice" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:SIQ\:SSS_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:SIQ\:SST_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:SIQ\:WS_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:SIQ\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:SIQ\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:SIQ\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:SIQ\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:SIQ\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:SIQ\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:SIQ\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:SIQ\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:SIQ\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:SIQ\:Poor_Quality = "64" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:SIQ\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:SIQ\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:Retrieval_Scheme = "3" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:Land_Rejected = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:Too_Close_To_Land_Rejected = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:Ice_Rejected = "10855" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:Missing_ECMWF_Rejected = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:Too_Few_Measurements_Rejected = "18084" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:Good_Quality_Grid_Points = "29636" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:Poor_Quality_Grid_Points = "4896" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:SQ\:Grid_Point_Type = "Sea" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:SQ\:SSS_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:SQ\:SST_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:SQ\:WS_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:SQ\:Good_Quality = "23293" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:SQ\:Good_Quality_Retrieved = "17816" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:SQ\:Good_Quality_Retrieved_Average_Sigma = "1.959542" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:SQ\:Good_Quality_Failed_Outside_Valid_Range = "81" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:SQ\:Good_Quality_Failed_Sigma_Too_High = "478" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:SQ\:Good_Quality_Failed_Poor_Fit = "5037" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:SQ\:Good_Quality_Failed_Marquardt = "4" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:SQ\:Good_Quality_Failed_Maxiter = "110" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:SQ\:Good_Quality_Failed_OOLUT = "555" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:SQ\:Poor_Quality = "2426" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:SQ\:Poor_Quality_Retrieved = "1661" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:SQ\:Poor_Quality_Retrieved_Average_Sigma = "2.933723" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:NCQ\:Grid_Point_Type = "Near_Coast" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:NCQ\:SSS_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:NCQ\:SST_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:NCQ\:WS_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:NCQ\:Good_Quality = "6343" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:NCQ\:Good_Quality_Retrieved = "3803" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:NCQ\:Good_Quality_Retrieved_Average_Sigma = "1.253443" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:NCQ\:Good_Quality_Failed_Outside_Valid_Range = "276" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:NCQ\:Good_Quality_Failed_Sigma_Too_High = "522" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:NCQ\:Good_Quality_Failed_Poor_Fit = "2247" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:NCQ\:Good_Quality_Failed_Marquardt = "152" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:NCQ\:Good_Quality_Failed_Maxiter = "411" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:NCQ\:Good_Quality_Failed_OOLUT = "773" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:NCQ\:Poor_Quality = "2470" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:NCQ\:Poor_Quality_Retrieved = "1367" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:NCQ\:Poor_Quality_Retrieved_Average_Sigma = "1.480500" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_0\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_0\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_0\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_0\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_0\:Good_Quality = "559" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_0\:Good_Quality_Retrieved = "131" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_0\:Good_Quality_Retrieved_Average_Sigma = "1.985529" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_0\:Good_Quality_Failed_Outside_Valid_Range = "183" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_0\:Good_Quality_Failed_Sigma_Too_High = "261" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_0\:Good_Quality_Failed_Poor_Fit = "325" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_0\:Good_Quality_Failed_Marquardt = "112" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_0\:Good_Quality_Failed_Maxiter = "130" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_0\:Good_Quality_Failed_OOLUT = "326" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_0\:Poor_Quality = "106" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_0\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_0\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_1\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_1\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_1\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_1\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_1\:Good_Quality = "486" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_1\:Good_Quality_Retrieved = "229" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_1\:Good_Quality_Retrieved_Average_Sigma = "2.167454" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_1\:Good_Quality_Failed_Outside_Valid_Range = "60" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_1\:Good_Quality_Failed_Sigma_Too_High = "82" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_1\:Good_Quality_Failed_Poor_Fit = "244" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_1\:Good_Quality_Failed_Marquardt = "30" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_1\:Good_Quality_Failed_Maxiter = "45" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_1\:Good_Quality_Failed_OOLUT = "135" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_1\:Poor_Quality = "233" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_1\:Poor_Quality_Retrieved = "13" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_1\:Poor_Quality_Retrieved_Average_Sigma = "4.597799" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_2\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_2\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_2\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_2\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_2\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_2\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_2\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_2\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_2\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_2\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_2\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_2\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_2\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_2\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_2\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_2\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_3\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_3\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_3\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_3\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_3\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_3\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_3\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_3\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_3\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_3\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_3\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_3\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_3\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_3\:Poor_Quality = "3" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_3\:Poor_Quality_Retrieved = "1" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_3\:Poor_Quality_Retrieved_Average_Sigma = "2.726585" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_4\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_4\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_4\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_4\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_4\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_4\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_4\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_4\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_4\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_4\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_4\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_4\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_4\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_4\:Poor_Quality = "233" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_4\:Poor_Quality_Retrieved = "182" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_4\:Poor_Quality_Retrieved_Average_Sigma = "3.945308" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_5\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_5\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_5\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_5\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_5\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_5\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_5\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_5\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_5\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_5\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_5\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_5\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_5\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_5\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_5\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_5\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_6\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_6\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_6\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_6\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_6\:Good_Quality = "16" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_6\:Good_Quality_Retrieved = "14" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_6\:Good_Quality_Retrieved_Average_Sigma = "1.307737" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_6\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_6\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_6\:Good_Quality_Failed_Poor_Fit = "2" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_6\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_6\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_6\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_6\:Poor_Quality = "22" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_6\:Poor_Quality_Retrieved = "19" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_6\:Poor_Quality_Retrieved_Average_Sigma = "1.902701" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_7\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_7\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_7\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_7\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_7\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_7\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_7\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_7\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_7\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_7\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_7\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_7\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_7\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_7\:Poor_Quality = "113" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_7\:Poor_Quality_Retrieved = "58" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_7\:Poor_Quality_Retrieved_Average_Sigma = "1.925949" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_8\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_8\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_8\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_8\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_8\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_8\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_8\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_8\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_8\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_8\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_8\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_8\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_8\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_8\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_8\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_8\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_9\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_9\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_9\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_9\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_9\:Good_Quality = "1485" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_9\:Good_Quality_Retrieved = "825" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_9\:Good_Quality_Retrieved_Average_Sigma = "2.191673" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_9\:Good_Quality_Failed_Outside_Valid_Range = "1" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_9\:Good_Quality_Failed_Sigma_Too_High = "54" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_9\:Good_Quality_Failed_Poor_Fit = "544" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_9\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_9\:Good_Quality_Failed_Maxiter = "247" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_9\:Good_Quality_Failed_OOLUT = "190" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_9\:Poor_Quality = "11" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_9\:Poor_Quality_Retrieved = "1" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_9\:Poor_Quality_Retrieved_Average_Sigma = "4.534814" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_10\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_10\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_10\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_10\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_10\:Good_Quality = "6940" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_10\:Good_Quality_Retrieved = "4685" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_10\:Good_Quality_Retrieved_Average_Sigma = "2.611991" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_10\:Good_Quality_Failed_Outside_Valid_Range = "102" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_10\:Good_Quality_Failed_Sigma_Too_High = "600" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_10\:Good_Quality_Failed_Poor_Fit = "1779" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_10\:Good_Quality_Failed_Marquardt = "14" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_10\:Good_Quality_Failed_Maxiter = "72" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_10\:Good_Quality_Failed_OOLUT = "603" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_10\:Poor_Quality = "508" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_10\:Poor_Quality_Retrieved = "218" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_10\:Poor_Quality_Retrieved_Average_Sigma = "4.334874" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_11\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_11\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_11\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_11\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_11\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_11\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_11\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_11\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_11\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_11\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_11\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_11\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_11\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_11\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_11\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_11\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_12\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_12\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_12\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_12\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_12\:Good_Quality = "232" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_12\:Good_Quality_Retrieved = "156" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_12\:Good_Quality_Retrieved_Average_Sigma = "1.521774" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_12\:Good_Quality_Failed_Outside_Valid_Range = "1" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_12\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_12\:Good_Quality_Failed_Poor_Fit = "70" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_12\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_12\:Good_Quality_Failed_Maxiter = "7" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_12\:Good_Quality_Failed_OOLUT = "17" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_12\:Poor_Quality = "55" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_12\:Poor_Quality_Retrieved = "42" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_12\:Poor_Quality_Retrieved_Average_Sigma = "2.482193" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_13\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_13\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_13\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_13\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_13\:Good_Quality = "11990" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_13\:Good_Quality_Retrieved = "9532" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_13\:Good_Quality_Retrieved_Average_Sigma = "2.064730" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_13\:Good_Quality_Failed_Outside_Valid_Range = "10" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_13\:Good_Quality_Failed_Sigma_Too_High = "3" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_13\:Good_Quality_Failed_Poor_Fit = "2454" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_13\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_13\:Good_Quality_Failed_Maxiter = "1" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_13\:Good_Quality_Failed_OOLUT = "42" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_13\:Poor_Quality = "997" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_13\:Poor_Quality_Retrieved = "857" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_13\:Poor_Quality_Retrieved_Average_Sigma = "3.092174" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_14\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_14\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_14\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_14\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_14\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_14\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_14\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_14\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_14\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_14\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_14\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_14\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_14\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_14\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_14\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_14\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_15\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_15\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_15\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_15\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_15\:Good_Quality = "830" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_15\:Good_Quality_Retrieved = "677" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_15\:Good_Quality_Retrieved_Average_Sigma = "1.047869" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_15\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_15\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_15\:Good_Quality_Failed_Poor_Fit = "153" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_15\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_15\:Good_Quality_Failed_Maxiter = "1" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_15\:Good_Quality_Failed_OOLUT = "4" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_15\:Poor_Quality = "1379" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_15\:Poor_Quality_Retrieved = "1092" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_15\:Poor_Quality_Retrieved_Average_Sigma = "1.087475" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_16\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_16\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_16\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_16\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_16\:Good_Quality = "7097" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_16\:Good_Quality_Retrieved = "5369" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_16\:Good_Quality_Retrieved_Average_Sigma = "0.787403" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_16\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_16\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_16\:Good_Quality_Failed_Poor_Fit = "1713" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_16\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_16\:Good_Quality_Failed_Maxiter = "18" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_16\:Good_Quality_Failed_OOLUT = "11" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_16\:Poor_Quality = "1043" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_16\:Poor_Quality_Retrieved = "450" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_16\:Poor_Quality_Retrieved_Average_Sigma = "1.581808" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_17\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_17\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_17\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_17\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_17\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_17\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_17\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_17\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_17\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_17\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_17\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_17\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_17\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_17\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_17\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_17\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_18\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_18\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_18\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_18\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_18\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_18\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_18\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_18\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_18\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_18\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_18\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_18\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_18\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_18\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_18\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_18\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_19\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_19\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_19\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_19\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_19\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_19\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_19\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_19\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_19\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_19\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_19\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_19\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_19\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_19\:Poor_Quality = "141" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_19\:Poor_Quality_Retrieved = "51" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_19\:Poor_Quality_Retrieved_Average_Sigma = "4.372903" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_20\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_20\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_20\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_20\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_20\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_20\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_20\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_20\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_20\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_20\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_20\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_20\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_20\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_20\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_20\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_20\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_21\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_21\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_21\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_21\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_21\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_21\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_21\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_21\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_21\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_21\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_21\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_21\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_21\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_21\:Poor_Quality = "8" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_21\:Poor_Quality_Retrieved = "5" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_21\:Poor_Quality_Retrieved_Average_Sigma = "2.769263" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_22\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_22\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_22\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_22\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_22\:Good_Quality = "1" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_22\:Good_Quality_Retrieved = "1" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_22\:Good_Quality_Retrieved_Average_Sigma = "2.597888" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_22\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_22\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_22\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_22\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_22\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_22\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_22\:Poor_Quality = "42" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_22\:Poor_Quality_Retrieved = "37" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_22\:Poor_Quality_Retrieved_Average_Sigma = "3.355307" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_23\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_23\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_23\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_23\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_23\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_23\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_23\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_23\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_23\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_23\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_23\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_23\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_23\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_23\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_23\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_23\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_24\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_24\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_24\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_24\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_24\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_24\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_24\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_24\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_24\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_24\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_24\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_24\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_24\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_24\:Poor_Quality = "2" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_24\:Poor_Quality_Retrieved = "2" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_24\:Poor_Quality_Retrieved_Average_Sigma = "2.113266" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_25\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_25\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_25\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_25\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_25\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_25\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_25\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_25\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_25\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_25\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_25\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_25\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_25\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_25\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_25\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_25\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_26\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_26\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_26\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_26\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_26\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_26\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_26\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_26\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_26\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_26\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_26\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_26\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_26\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_26\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_26\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_26\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:SIQ\:Grid_Point_Type = "Sea_Ice" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:SIQ\:SSS_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:SIQ\:SST_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:SIQ\:WS_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:SIQ\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:SIQ\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:SIQ\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:SIQ\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:SIQ\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:SIQ\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:SIQ\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:SIQ\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:SIQ\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:SIQ\:Poor_Quality = "64" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:SIQ\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:SIQ\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:Retrieval_Scheme = "4" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:Land_Rejected = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:Too_Close_To_Land_Rejected = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:Ice_Rejected = "10855" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:Missing_ECMWF_Rejected = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:Too_Few_Measurements_Rejected = "18084" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:Good_Quality_Grid_Points = "29899" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:Poor_Quality_Grid_Points = "4633" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:SQ\:Grid_Point_Type = "Sea" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:SQ\:SSS_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:SQ\:SST_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:SQ\:WS_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:SQ\:Good_Quality = "23293" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:SQ\:Good_Quality_Retrieved = "21547" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:SQ\:Good_Quality_Retrieved_Average_Sigma = "0.736739" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:SQ\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:SQ\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:SQ\:Good_Quality_Failed_Poor_Fit = "1746" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:SQ\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:SQ\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:SQ\:Good_Quality_Failed_OOLUT = "1638" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:SQ\:Poor_Quality = "2426" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:SQ\:Poor_Quality_Retrieved = "1988" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:SQ\:Poor_Quality_Retrieved_Average_Sigma = "1.498341" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:NCQ\:Grid_Point_Type = "Near_Coast" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:NCQ\:SSS_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:NCQ\:SST_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:NCQ\:WS_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:NCQ\:Good_Quality = "6606" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:NCQ\:Good_Quality_Retrieved = "5264" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:NCQ\:Good_Quality_Retrieved_Average_Sigma = "0.828990" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:NCQ\:Good_Quality_Failed_Outside_Valid_Range = "254" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:NCQ\:Good_Quality_Failed_Sigma_Too_High = "32" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:NCQ\:Good_Quality_Failed_Poor_Fit = "1330" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:NCQ\:Good_Quality_Failed_Marquardt = "8" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:NCQ\:Good_Quality_Failed_Maxiter = "2" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:NCQ\:Good_Quality_Failed_OOLUT = "927" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:NCQ\:Poor_Quality = "2207" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:NCQ\:Poor_Quality_Retrieved = "1429" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:NCQ\:Poor_Quality_Retrieved_Average_Sigma = "1.448753" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_0\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_0\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_0\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_0\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_0\:Good_Quality = "559" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_0\:Good_Quality_Retrieved = "358" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_0\:Good_Quality_Retrieved_Average_Sigma = "0.674638" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_0\:Good_Quality_Failed_Outside_Valid_Range = "30" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_0\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_0\:Good_Quality_Failed_Poor_Fit = "190" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_0\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_0\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_0\:Good_Quality_Failed_OOLUT = "201" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_0\:Poor_Quality = "106" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_0\:Poor_Quality_Retrieved = "29" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_0\:Poor_Quality_Retrieved_Average_Sigma = "1.338563" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_1\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_1\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_1\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_1\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_1\:Good_Quality = "486" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_1\:Good_Quality_Retrieved = "385" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_1\:Good_Quality_Retrieved_Average_Sigma = "0.616946" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_1\:Good_Quality_Failed_Outside_Valid_Range = "4" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_1\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_1\:Good_Quality_Failed_Poor_Fit = "101" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_1\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_1\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_1\:Good_Quality_Failed_OOLUT = "101" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_1\:Poor_Quality = "233" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_1\:Poor_Quality_Retrieved = "136" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_1\:Poor_Quality_Retrieved_Average_Sigma = "1.539670" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_2\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_2\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_2\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_2\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_2\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_2\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_2\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_2\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_2\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_2\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_2\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_2\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_2\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_2\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_2\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_2\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_3\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_3\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_3\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_3\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_3\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_3\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_3\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_3\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_3\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_3\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_3\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_3\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_3\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_3\:Poor_Quality = "3" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_3\:Poor_Quality_Retrieved = "1" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_3\:Poor_Quality_Retrieved_Average_Sigma = "2.143224" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_4\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_4\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_4\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_4\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_4\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_4\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_4\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_4\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_4\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_4\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_4\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_4\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_4\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_4\:Poor_Quality = "233" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_4\:Poor_Quality_Retrieved = "187" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_4\:Poor_Quality_Retrieved_Average_Sigma = "1.582498" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_5\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_5\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_5\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_5\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_5\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_5\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_5\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_5\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_5\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_5\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_5\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_5\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_5\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_5\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_5\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_5\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_6\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_6\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_6\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_6\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_6\:Good_Quality = "16" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_6\:Good_Quality_Retrieved = "15" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_6\:Good_Quality_Retrieved_Average_Sigma = "1.357438" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_6\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_6\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_6\:Good_Quality_Failed_Poor_Fit = "1" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_6\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_6\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_6\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_6\:Poor_Quality = "22" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_6\:Poor_Quality_Retrieved = "19" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_6\:Poor_Quality_Retrieved_Average_Sigma = "2.030221" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_7\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_7\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_7\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_7\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_7\:Good_Quality = "28" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_7\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_7\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_7\:Good_Quality_Failed_Outside_Valid_Range = "19" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_7\:Good_Quality_Failed_Sigma_Too_High = "4" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_7\:Good_Quality_Failed_Poor_Fit = "28" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_7\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_7\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_7\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_7\:Poor_Quality = "85" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_7\:Poor_Quality_Retrieved = "53" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_7\:Poor_Quality_Retrieved_Average_Sigma = "1.845069" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_8\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_8\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_8\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_8\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_8\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_8\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_8\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_8\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_8\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_8\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_8\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_8\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_8\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_8\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_8\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_8\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_9\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_9\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_9\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_9\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_9\:Good_Quality = "1485" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_9\:Good_Quality_Retrieved = "1275" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_9\:Good_Quality_Retrieved_Average_Sigma = "0.643317" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_9\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_9\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_9\:Good_Quality_Failed_Poor_Fit = "210" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_9\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_9\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_9\:Good_Quality_Failed_OOLUT = "210" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_9\:Poor_Quality = "11" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_9\:Poor_Quality_Retrieved = "6" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_9\:Poor_Quality_Retrieved_Average_Sigma = "1.393877" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_10\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_10\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_10\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_10\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_10\:Good_Quality = "6940" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_10\:Good_Quality_Retrieved = "6223" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_10\:Good_Quality_Retrieved_Average_Sigma = "0.743647" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_10\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_10\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_10\:Good_Quality_Failed_Poor_Fit = "717" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_10\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_10\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_10\:Good_Quality_Failed_OOLUT = "717" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_10\:Poor_Quality = "508" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_10\:Poor_Quality_Retrieved = "387" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_10\:Poor_Quality_Retrieved_Average_Sigma = "1.451606" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_11\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_11\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_11\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_11\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_11\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_11\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_11\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_11\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_11\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_11\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_11\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_11\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_11\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_11\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_11\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_11\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_12\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_12\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_12\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_12\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_12\:Good_Quality = "232" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_12\:Good_Quality_Retrieved = "213" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_12\:Good_Quality_Retrieved_Average_Sigma = "0.741777" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_12\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_12\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_12\:Good_Quality_Failed_Poor_Fit = "19" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_12\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_12\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_12\:Good_Quality_Failed_OOLUT = "17" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_12\:Poor_Quality = "55" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_12\:Poor_Quality_Retrieved = "42" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_12\:Poor_Quality_Retrieved_Average_Sigma = "2.121626" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_13\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_13\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_13\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_13\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_13\:Good_Quality = "11990" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_13\:Good_Quality_Retrieved = "11136" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_13\:Good_Quality_Retrieved_Average_Sigma = "0.731001" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_13\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_13\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_13\:Good_Quality_Failed_Poor_Fit = "854" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_13\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_13\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_13\:Good_Quality_Failed_OOLUT = "813" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_13\:Poor_Quality = "997" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_13\:Poor_Quality_Retrieved = "847" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_13\:Poor_Quality_Retrieved_Average_Sigma = "1.560844" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_14\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_14\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_14\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_14\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_14\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_14\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_14\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_14\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_14\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_14\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_14\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_14\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_14\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_14\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_14\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_14\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_15\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_15\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_15\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_15\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_15\:Good_Quality = "830" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_15\:Good_Quality_Retrieved = "722" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_15\:Good_Quality_Retrieved_Average_Sigma = "1.117939" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_15\:Good_Quality_Failed_Outside_Valid_Range = "1" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_15\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_15\:Good_Quality_Failed_Poor_Fit = "107" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_15\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_15\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_15\:Good_Quality_Failed_OOLUT = "39" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_15\:Poor_Quality = "1379" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_15\:Poor_Quality_Retrieved = "1079" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_15\:Poor_Quality_Retrieved_Average_Sigma = "1.235114" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_16\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_16\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_16\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_16\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_16\:Good_Quality = "7332" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_16\:Good_Quality_Retrieved = "6483" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_16\:Good_Quality_Retrieved_Average_Sigma = "0.799682" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_16\:Good_Quality_Failed_Outside_Valid_Range = "200" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_16\:Good_Quality_Failed_Sigma_Too_High = "28" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_16\:Good_Quality_Failed_Poor_Fit = "849" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_16\:Good_Quality_Failed_Marquardt = "8" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_16\:Good_Quality_Failed_Maxiter = "2" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_16\:Good_Quality_Failed_OOLUT = "467" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_16\:Poor_Quality = "808" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_16\:Poor_Quality_Retrieved = "463" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_16\:Poor_Quality_Retrieved_Average_Sigma = "1.640629" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_17\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_17\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_17\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_17\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_17\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_17\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_17\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_17\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_17\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_17\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_17\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_17\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_17\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_17\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_17\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_17\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_18\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_18\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_18\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_18\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_18\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_18\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_18\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_18\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_18\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_18\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_18\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_18\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_18\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_18\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_18\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_18\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_19\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_19\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_19\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_19\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_19\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_19\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_19\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_19\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_19\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_19\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_19\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_19\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_19\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_19\:Poor_Quality = "141" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_19\:Poor_Quality_Retrieved = "127" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_19\:Poor_Quality_Retrieved_Average_Sigma = "1.663481" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_20\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_20\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_20\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_20\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_20\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_20\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_20\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_20\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_20\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_20\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_20\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_20\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_20\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_20\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_20\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_20\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_21\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_21\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_21\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_21\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_21\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_21\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_21\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_21\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_21\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_21\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_21\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_21\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_21\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_21\:Poor_Quality = "8" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_21\:Poor_Quality_Retrieved = "5" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_21\:Poor_Quality_Retrieved_Average_Sigma = "2.440643" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_22\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_22\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_22\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_22\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_22\:Good_Quality = "1" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_22\:Good_Quality_Retrieved = "1" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_22\:Good_Quality_Retrieved_Average_Sigma = "1.041794" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_22\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_22\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_22\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_22\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_22\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_22\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_22\:Poor_Quality = "42" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_22\:Poor_Quality_Retrieved = "36" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_22\:Poor_Quality_Retrieved_Average_Sigma = "1.924485" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_23\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_23\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_23\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_23\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_23\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_23\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_23\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_23\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_23\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_23\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_23\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_23\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_23\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_23\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_23\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_23\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_24\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_24\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_24\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_24\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_24\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_24\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_24\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_24\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_24\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_24\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_24\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_24\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_24\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_24\:Poor_Quality = "2" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_24\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_24\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_25\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_25\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_25\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_25\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_25\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_25\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_25\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_25\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_25\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_25\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_25\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_25\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_25\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_25\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_25\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_25\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_26\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_26\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_26\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_26\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_26\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_26\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_26\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_26\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_26\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_26\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_26\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_26\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_26\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_26\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_26\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_26\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:SIQ\:Grid_Point_Type = "Sea_Ice" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:SIQ\:SSS_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:SIQ\:SST_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:SIQ\:WS_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:SIQ\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:SIQ\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:SIQ\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:SIQ\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:SIQ\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:SIQ\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:SIQ\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:SIQ\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:SIQ\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:SIQ\:Poor_Quality = "64" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:SIQ\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:SIQ\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_0\:Retrieved_Parameter_0\:name = "SSS" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_0\:Retrieved_Parameter_0\:unit = "Practical Salinity Unit (PSU)" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_0\:Retrieved_Parameter_0\:description = "Surface salinity of the sea at gridpoint" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_0\:Retrieved_Parameter_1\:name = "SST" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_0\:Retrieved_Parameter_1\:unit = "Kelvin" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_0\:Retrieved_Parameter_1\:description = "Surface temperature of the sea at gridpoint" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_0\:Retrieved_Parameter_2\:name = "UN10" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_0\:Retrieved_Parameter_2\:unit = "m.s-1" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_0\:Retrieved_Parameter_2\:description = "U component of neutral wind 10m above surface" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_0\:Retrieved_Parameter_3\:name = "VN10" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_0\:Retrieved_Parameter_3\:unit = "m.s-1" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_0\:Retrieved_Parameter_3\:description = "V component of neutral wind 10m above surface" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_0\:Retrieved_Parameter_4\:name = "tec" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_0\:Retrieved_Parameter_4\:unit = "tecu" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_0\:Retrieved_Parameter_4\:description = "Total Electronic Content of the ionosphere below SMOS" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_0\:Retrieved_Parameter_5\:name = "not used" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_0\:Retrieved_Parameter_5\:unit = "none" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_0\:Retrieved_Parameter_5\:description = "no parameter defined" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_0\:Retrieved_Parameter_6\:name = "not used" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_0\:Retrieved_Parameter_6\:unit = "none" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_0\:Retrieved_Parameter_6\:description = "no parameter defined" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_0\:Retrieved_Parameter_7\:name = "not used" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_0\:Retrieved_Parameter_7\:unit = "none" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_0\:Retrieved_Parameter_7\:description = "no parameter defined" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_0\:Retrieved_Parameter_8\:name = "not used" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_0\:Retrieved_Parameter_8\:unit = "none" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_0\:Retrieved_Parameter_8\:description = "no parameter defined" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_0\:Retrieved_Parameter_9\:name = "not used" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_0\:Retrieved_Parameter_9\:unit = "none" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_0\:Retrieved_Parameter_9\:description = "no parameter defined" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_1\:Retrieved_Parameter_0\:name = "SSS" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_1\:Retrieved_Parameter_0\:unit = "Practical Salinity Unit (PSU)" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_1\:Retrieved_Parameter_0\:description = "Surface salinity of the sea at gridpoint" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_1\:Retrieved_Parameter_1\:name = "SST" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_1\:Retrieved_Parameter_1\:unit = "Kelvin" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_1\:Retrieved_Parameter_1\:description = "Surface temperature of the sea at gridpoint" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_1\:Retrieved_Parameter_2\:name = "UN10" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_1\:Retrieved_Parameter_2\:unit = "m.s-1" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_1\:Retrieved_Parameter_2\:description = "U component of neutral wind 10m above surface" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_1\:Retrieved_Parameter_3\:name = "VN10" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_1\:Retrieved_Parameter_3\:unit = "m.s-1" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_1\:Retrieved_Parameter_3\:description = "V component of neutral wind 10m above surface" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_1\:Retrieved_Parameter_4\:name = "tec" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_1\:Retrieved_Parameter_4\:unit = "tecu" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_1\:Retrieved_Parameter_4\:description = "Total Electronic Content of the ionosphere below SMOS" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_1\:Retrieved_Parameter_5\:name = "not used" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_1\:Retrieved_Parameter_5\:unit = "none" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_1\:Retrieved_Parameter_5\:description = "no parameter defined" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_1\:Retrieved_Parameter_6\:name = "not used" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_1\:Retrieved_Parameter_6\:unit = "none" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_1\:Retrieved_Parameter_6\:description = "no parameter defined" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_1\:Retrieved_Parameter_7\:name = "not used" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_1\:Retrieved_Parameter_7\:unit = "none" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_1\:Retrieved_Parameter_7\:description = "no parameter defined" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_1\:Retrieved_Parameter_8\:name = "not used" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_1\:Retrieved_Parameter_8\:unit = "none" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_1\:Retrieved_Parameter_8\:description = "no parameter defined" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_1\:Retrieved_Parameter_9\:name = "not used" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_1\:Retrieved_Parameter_9\:unit = "none" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_1\:Retrieved_Parameter_9\:description = "no parameter defined" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_2\:Retrieved_Parameter_0\:name = "SSS" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_2\:Retrieved_Parameter_0\:unit = "Practical Salinity Unit (PSU)" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_2\:Retrieved_Parameter_0\:description = "Surface salinity of the sea at gridpoint" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_2\:Retrieved_Parameter_1\:name = "SST" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_2\:Retrieved_Parameter_1\:unit = "Kelvin" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_2\:Retrieved_Parameter_1\:description = "Surface temperature of the sea at gridpoint" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_2\:Retrieved_Parameter_2\:name = "UN10" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_2\:Retrieved_Parameter_2\:unit = "m.s-1" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_2\:Retrieved_Parameter_2\:description = "U component of neutral wind 10m above surface" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_2\:Retrieved_Parameter_3\:name = "VN10" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_2\:Retrieved_Parameter_3\:unit = "m.s-1" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_2\:Retrieved_Parameter_3\:description = "V component of neutral wind 10m above surface" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_2\:Retrieved_Parameter_4\:name = "tec" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_2\:Retrieved_Parameter_4\:unit = "tecu" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_2\:Retrieved_Parameter_4\:description = "Total Electronic Content of the ionosphere below SMOS" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_2\:Retrieved_Parameter_5\:name = "not used" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_2\:Retrieved_Parameter_5\:unit = "none" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_2\:Retrieved_Parameter_5\:description = "no parameter defined" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_2\:Retrieved_Parameter_6\:name = "not used" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_2\:Retrieved_Parameter_6\:unit = "none" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_2\:Retrieved_Parameter_6\:description = "no parameter defined" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_2\:Retrieved_Parameter_7\:name = "not used" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_2\:Retrieved_Parameter_7\:unit = "none" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_2\:Retrieved_Parameter_7\:description = "no parameter defined" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_2\:Retrieved_Parameter_8\:name = "not used" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_2\:Retrieved_Parameter_8\:unit = "none" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_2\:Retrieved_Parameter_8\:description = "no parameter defined" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_2\:Retrieved_Parameter_9\:name = "not used" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_2\:Retrieved_Parameter_9\:unit = "none" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_2\:Retrieved_Parameter_9\:description = "no parameter defined" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_3\:Retrieved_Parameter_0\:name = "Acard" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_3\:Retrieved_Parameter_0\:unit = "dl" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_3\:Retrieved_Parameter_0\:description = "Acard coefficient for cardioid model" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_3\:Retrieved_Parameter_1\:name = "SST" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_3\:Retrieved_Parameter_1\:unit = "Kelvin" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_3\:Retrieved_Parameter_1\:description = "Surface temperature of the sea at gridpoint" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_3\:Retrieved_Parameter_2\:name = "not used" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_3\:Retrieved_Parameter_2\:unit = "none" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_3\:Retrieved_Parameter_2\:description = "no parameter defined" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_3\:Retrieved_Parameter_3\:name = "not used" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_3\:Retrieved_Parameter_3\:unit = "none" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_3\:Retrieved_Parameter_3\:description = "no parameter defined" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_3\:Retrieved_Parameter_4\:name = "not used" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_3\:Retrieved_Parameter_4\:unit = "none" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_3\:Retrieved_Parameter_4\:description = "no parameter defined" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_3\:Retrieved_Parameter_5\:name = "not used" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_3\:Retrieved_Parameter_5\:unit = "none" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_3\:Retrieved_Parameter_5\:description = "no parameter defined" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_3\:Retrieved_Parameter_6\:name = "not used" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_3\:Retrieved_Parameter_6\:unit = "none" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_3\:Retrieved_Parameter_6\:description = "no parameter defined" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_3\:Retrieved_Parameter_7\:name = "not used" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_3\:Retrieved_Parameter_7\:unit = "none" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_3\:Retrieved_Parameter_7\:description = "no parameter defined" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_3\:Retrieved_Parameter_8\:name = "not used" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_3\:Retrieved_Parameter_8\:unit = "none" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_3\:Retrieved_Parameter_8\:description = "no parameter defined" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_3\:Retrieved_Parameter_9\:name = "not used" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_3\:Retrieved_Parameter_9\:unit = "none" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_3\:Retrieved_Parameter_9\:description = "no parameter defined" ;
		string :VH\:SPH\:MI\:SPH_Descriptor = "MIR_OSUDP2_SPH" ;
		string :VH\:SPH\:MI\:Checksum = "0186172426" ;
		string :VH\:SPH\:MI\:Header_Schema = "HDR_SM_XXXX_MIR_OSUDP2_0400.xsd" ;
		string :VH\:SPH\:MI\:Datablock_Schema = "DBL_SM_XXXX_MIR_OSUDP2_0401.binXschema.xml" ;
		string :VH\:SPH\:MI\:Header_Size = "168617" ;
		string :VH\:SPH\:MI\:Datablock_Size = "00017615474" ;
		string :VH\:SPH\:MI\:HW_Identifier = "0002" ;
		string :VH\:SPH\:MI\:TI\:Precise_Validity_Start = "UTC=2021-06-30T21:59:10.071954" ;
		string :VH\:SPH\:MI\:TI\:Precise_Validity_Stop = "UTC=2021-06-30T22:52:30.511865" ;
		string :VH\:SPH\:MI\:TI\:Abs_Orbit_Start = "+61281" ;
		string :VH\:SPH\:MI\:TI\:Start_Time_ANX_T = "4283.930491" ;
		string :VH\:SPH\:MI\:TI\:Abs_Orbit_Stop = "+61282" ;
		string :VH\:SPH\:MI\:TI\:Stop_Time_ANX_T = "1479.892790" ;
		string :VH\:SPH\:MI\:TI\:UTC_at_ANX = "UTC=2021-06-30T20:47:46.141463" ;
		string :VH\:SPH\:MI\:TI\:Long_at_ANX = "+138.381497" ;
		string :VH\:SPH\:MI\:TI\:Ascending_Flag = "A" ;
		string :VH\:SPH\:MI\:TI\:Polarisation_Flag = "F" ;
		string :VH\:SPH\:LODS\:Data_Set_0\:DS_Name = "SSS_SWATH" ;
		string :VH\:SPH\:LODS\:Data_Set_0\:DS_Type = "M" ;
		string :VH\:SPH\:LODS\:Data_Set_0\:DS_Size = "0017615474" ;
		string :VH\:SPH\:LODS\:Data_Set_0\:DS_Offset = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_0\:Num_DSR = "0000092713" ;
		string :VH\:SPH\:LODS\:Data_Set_0\:DSR_Size = "00000190" ;
		string :VH\:SPH\:LODS\:Data_Set_0\:Byte_Order = "0123" ;
		string :VH\:SPH\:LODS\:Data_Set_1\:DS_Name = "L1C_OS_FILE" ;
		string :VH\:SPH\:LODS\:Data_Set_1\:DS_Type = "R" ;
		string :VH\:SPH\:LODS\:Data_Set_1\:DS_Size = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_1\:DS_Offset = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_1\:Ref_Filename = "SM_OPER_MIR_SCSF1C_20210630T215911_20210630T225230_724_001_1" ;
		string :VH\:SPH\:LODS\:Data_Set_1\:Num_DSR = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_1\:DSR_Size = "00000000" ;
		string :VH\:SPH\:LODS\:Data_Set_1\:Byte_Order = "0000" ;
		string :VH\:SPH\:LODS\:Data_Set_2\:DS_Name = "DGG_FILE" ;
		string :VH\:SPH\:LODS\:Data_Set_2\:DS_Type = "R" ;
		string :VH\:SPH\:LODS\:Data_Set_2\:DS_Size = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_2\:DS_Offset = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_2\:Ref_Filename = "SM_OPER_AUX_DGG____20050101T000000_20500101T000000_300_003_3" ;
		string :VH\:SPH\:LODS\:Data_Set_2\:Num_DSR = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_2\:DSR_Size = "00000000" ;
		string :VH\:SPH\:LODS\:Data_Set_2\:Byte_Order = "0000" ;
		string :VH\:SPH\:LODS\:Data_Set_3\:DS_Name = "IERS_BULLETIN_B_FILE" ;
		string :VH\:SPH\:LODS\:Data_Set_3\:DS_Type = "R" ;
		string :VH\:SPH\:LODS\:Data_Set_3\:DS_Size = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_3\:DS_Offset = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_3\:Ref_Filename = "SM_OPER_AUX_BULL_B_20210402T000000_20500101T000000_120_001_3" ;
		string :VH\:SPH\:LODS\:Data_Set_3\:Num_DSR = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_3\:DSR_Size = "00000000" ;
		string :VH\:SPH\:LODS\:Data_Set_3\:Byte_Order = "0000" ;
		string :VH\:SPH\:LODS\:Data_Set_4\:DS_Name = "BESTFITPLANE_FILE" ;
		string :VH\:SPH\:LODS\:Data_Set_4\:DS_Type = "R" ;
		string :VH\:SPH\:LODS\:Data_Set_4\:DS_Size = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_4\:DS_Offset = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_4\:Ref_Filename = "SM_OPER_AUX_BFP____20050101T000000_20500101T000000_340_004_3" ;
		string :VH\:SPH\:LODS\:Data_Set_4\:Num_DSR = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_4\:DSR_Size = "00000000" ;
		string :VH\:SPH\:LODS\:Data_Set_4\:Byte_Order = "0000" ;
		string :VH\:SPH\:LODS\:Data_Set_5\:DS_Name = "MISPOINTING_FILE" ;
		string :VH\:SPH\:LODS\:Data_Set_5\:DS_Type = "R" ;
		string :VH\:SPH\:LODS\:Data_Set_5\:DS_Size = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_5\:DS_Offset = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_5\:Ref_Filename = "SM_OPER_AUX_MISP___20050101T000000_20500101T000000_300_004_3" ;
		string :VH\:SPH\:LODS\:Data_Set_5\:Num_DSR = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_5\:DSR_Size = "00000000" ;
		string :VH\:SPH\:LODS\:Data_Set_5\:Byte_Order = "0000" ;
		string :VH\:SPH\:LODS\:Data_Set_6\:DS_Name = "ECMWF_FILE" ;
		string :VH\:SPH\:LODS\:Data_Set_6\:DS_Type = "R" ;
		string :VH\:SPH\:LODS\:Data_Set_6\:DS_Size = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_6\:DS_Offset = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_6\:Ref_Filename = "SM_OPER_AUX_ECMWF__20210630T215902_20210630T230542_318_001_3" ;
		string :VH\:SPH\:LODS\:Data_Set_6\:Num_DSR = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_6\:DSR_Size = "00000000" ;
		string :VH\:SPH\:LODS\:Data_Set_6\:Byte_Order = "0000" ;
		string :VH\:SPH\:LODS\:Data_Set_7\:DS_Name = "FLAT_SEA_FILE" ;
		string :VH\:SPH\:LODS\:Data_Set_7\:DS_Type = "R" ;
		string :VH\:SPH\:LODS\:Data_Set_7\:DS_Size = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_7\:DS_Offset = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_7\:Ref_Filename = "SM_OPER_AUX_FLTSEA_20050101T000000_20500101T000000_001_012_3" ;
		string :VH\:SPH\:LODS\:Data_Set_7\:Num_DSR = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_7\:DSR_Size = "00000000" ;
		string :VH\:SPH\:LODS\:Data_Set_7\:Byte_Order = "0000" ;
		string :VH\:SPH\:LODS\:Data_Set_8\:DS_Name = "ROUGHNESS_IPSL_FILE" ;
		string :VH\:SPH\:LODS\:Data_Set_8\:DS_Type = "R" ;
		string :VH\:SPH\:LODS\:Data_Set_8\:DS_Size = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_8\:DS_Offset = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_8\:Ref_Filename = "SM_OPER_AUX_RGHNS1_20050101T000000_20500101T000000_001_016_3" ;
		string :VH\:SPH\:LODS\:Data_Set_8\:Num_DSR = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_8\:DSR_Size = "00000000" ;
		string :VH\:SPH\:LODS\:Data_Set_8\:Byte_Order = "0000" ;
		string :VH\:SPH\:LODS\:Data_Set_9\:DS_Name = "ROUGHNESS_IFREMER_FILE" ;
		string :VH\:SPH\:LODS\:Data_Set_9\:DS_Type = "R" ;
		string :VH\:SPH\:LODS\:Data_Set_9\:DS_Size = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_9\:DS_Offset = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_9\:Ref_Filename = "SM_OPER_AUX_RGHNS2_20050101T000000_20500101T000000_001_013_3" ;
		string :VH\:SPH\:LODS\:Data_Set_9\:Num_DSR = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_9\:DSR_Size = "00000000" ;
		string :VH\:SPH\:LODS\:Data_Set_9\:Byte_Order = "0000" ;
		string :VH\:SPH\:LODS\:Data_Set_10\:DS_Name = "ROUGHNESS_ICM_CSIC_FILE" ;
		string :VH\:SPH\:LODS\:Data_Set_10\:DS_Type = "R" ;
		string :VH\:SPH\:LODS\:Data_Set_10\:DS_Size = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_10\:DS_Offset = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_10\:Ref_Filename = "SM_OPER_AUX_RGHNS3_20050101T000000_20500101T000000_001_016_3" ;
		string :VH\:SPH\:LODS\:Data_Set_10\:Num_DSR = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_10\:DSR_Size = "00000000" ;
		string :VH\:SPH\:LODS\:Data_Set_10\:Byte_Order = "0000" ;
		string :VH\:SPH\:LODS\:Data_Set_11\:DS_Name = "GALAXY_OS_FILE" ;
		string :VH\:SPH\:LODS\:Data_Set_11\:DS_Type = "R" ;
		string :VH\:SPH\:LODS\:Data_Set_11\:DS_Size = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_11\:DS_Offset = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_11\:Ref_Filename = "SM_OPER_AUX_GAL_OS_20050101T000000_20500101T000000_001_011_3" ;
		string :VH\:SPH\:LODS\:Data_Set_11\:Num_DSR = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_11\:DSR_Size = "00000000" ;
		string :VH\:SPH\:LODS\:Data_Set_11\:Byte_Order = "0000" ;
		string :VH\:SPH\:LODS\:Data_Set_12\:DS_Name = "GALAXY_2OS_FILE" ;
		string :VH\:SPH\:LODS\:Data_Set_12\:DS_Type = "R" ;
		string :VH\:SPH\:LODS\:Data_Set_12\:DS_Size = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_12\:DS_Offset = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_12\:Ref_Filename = "SM_OPER_AUX_GAL2OS_20050101T000000_20500101T000000_001_016_3" ;
		string :VH\:SPH\:LODS\:Data_Set_12\:Num_DSR = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_12\:DSR_Size = "00000000" ;
		string :VH\:SPH\:LODS\:Data_Set_12\:Byte_Order = "0000" ;
		string :VH\:SPH\:LODS\:Data_Set_13\:DS_Name = "SUNGLINT_FILE" ;
		string :VH\:SPH\:LODS\:Data_Set_13\:DS_Type = "R" ;
		string :VH\:SPH\:LODS\:Data_Set_13\:DS_Size = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_13\:DS_Offset = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_13\:Ref_Filename = "SM_OPER_AUX_SGLINT_20050101T000000_20500101T000000_001_012_3" ;
		string :VH\:SPH\:LODS\:Data_Set_13\:Num_DSR = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_13\:DSR_Size = "00000000" ;
		string :VH\:SPH\:LODS\:Data_Set_13\:Byte_Order = "0000" ;
		string :VH\:SPH\:LODS\:Data_Set_14\:DS_Name = "ATMOS_FILE" ;
		string :VH\:SPH\:LODS\:Data_Set_14\:DS_Type = "R" ;
		string :VH\:SPH\:LODS\:Data_Set_14\:DS_Size = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_14\:DS_Offset = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_14\:Ref_Filename = "SM_OPER_AUX_ATMOS__20050101T000000_20500101T000000_001_010_3" ;
		string :VH\:SPH\:LODS\:Data_Set_14\:Num_DSR = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_14\:DSR_Size = "00000000" ;
		string :VH\:SPH\:LODS\:Data_Set_14\:Byte_Order = "0000" ;
		string :VH\:SPH\:LODS\:Data_Set_15\:DS_Name = "DISTAN_FILE" ;
		string :VH\:SPH\:LODS\:Data_Set_15\:DS_Type = "R" ;
		string :VH\:SPH\:LODS\:Data_Set_15\:DS_Size = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_15\:DS_Offset = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_15\:Ref_Filename = "SM_OPER_AUX_DISTAN_20050101T000000_20500101T000000_001_011_3" ;
		string :VH\:SPH\:LODS\:Data_Set_15\:Num_DSR = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_15\:DSR_Size = "00000000" ;
		string :VH\:SPH\:LODS\:Data_Set_15\:Byte_Order = "0000" ;
		string :VH\:SPH\:LODS\:Data_Set_16\:DS_Name = "CLIMATOLOGY_SSS_FILE" ;
		string :VH\:SPH\:LODS\:Data_Set_16\:DS_Type = "R" ;
		string :VH\:SPH\:LODS\:Data_Set_16\:DS_Size = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_16\:DS_Offset = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_16\:Ref_Filename = "SM_OPER_AUX_SSS____20050101T000000_20500101T000000_001_014_3" ;
		string :VH\:SPH\:LODS\:Data_Set_16\:Num_DSR = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_16\:DSR_Size = "00000000" ;
		string :VH\:SPH\:LODS\:Data_Set_16\:Byte_Order = "0000" ;
		string :VH\:SPH\:LODS\:Data_Set_17\:DS_Name = "CLIMATOLOGY_SSSCLI_FILE" ;
		string :VH\:SPH\:LODS\:Data_Set_17\:DS_Type = "R" ;
		string :VH\:SPH\:LODS\:Data_Set_17\:DS_Size = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_17\:DS_Offset = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_17\:Ref_Filename = "SM_OPER_AUX_SSSCLI_20050101T000000_20500101T000000_001_002_3" ;
		string :VH\:SPH\:LODS\:Data_Set_17\:Num_DSR = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_17\:DSR_Size = "00000000" ;
		string :VH\:SPH\:LODS\:Data_Set_17\:Byte_Order = "0000" ;
		string :VH\:SPH\:LODS\:Data_Set_18\:DS_Name = "OCEAN_SALINITY_CONFIG_FILE" ;
		string :VH\:SPH\:LODS\:Data_Set_18\:DS_Type = "R" ;
		string :VH\:SPH\:LODS\:Data_Set_18\:DS_Size = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_18\:DS_Offset = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_18\:Ref_Filename = "SM_OPER_AUX_CNFOSF_20050101T000000_20500101T000000_001_032_3" ;
		string :VH\:SPH\:LODS\:Data_Set_18\:Num_DSR = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_18\:DSR_Size = "00000000" ;
		string :VH\:SPH\:LODS\:Data_Set_18\:Byte_Order = "0000" ;
		string :VH\:SPH\:LODS\:Data_Set_19\:DS_Name = "OTT1F_FILE" ;
		string :VH\:SPH\:LODS\:Data_Set_19\:DS_Type = "R" ;
		string :VH\:SPH\:LODS\:Data_Set_19\:DS_Size = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_19\:DS_Offset = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_19\:Ref_Filename = "SM_OPER_AUX_OTT1F__20210624T082406_20500101T000000_700_001_1" ;
		string :VH\:SPH\:LODS\:Data_Set_19\:Num_DSR = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_19\:DSR_Size = "00000000" ;
		string :VH\:SPH\:LODS\:Data_Set_19\:Byte_Order = "0000" ;
		string :VH\:SPH\:LODS\:Data_Set_20\:DS_Name = "OTT2F_FILE" ;
		string :VH\:SPH\:LODS\:Data_Set_20\:DS_Type = "R" ;
		string :VH\:SPH\:LODS\:Data_Set_20\:DS_Size = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_20\:DS_Offset = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_20\:Ref_Filename = "SM_OPER_AUX_OTT2F__20210624T082406_20500101T000000_700_001_1" ;
		string :VH\:SPH\:LODS\:Data_Set_20\:Num_DSR = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_20\:DSR_Size = "00000000" ;
		string :VH\:SPH\:LODS\:Data_Set_20\:Byte_Order = "0000" ;
		string :VH\:SPH\:LODS\:Data_Set_21\:DS_Name = "OTT3F_FILE" ;
		string :VH\:SPH\:LODS\:Data_Set_21\:DS_Type = "R" ;
		string :VH\:SPH\:LODS\:Data_Set_21\:DS_Size = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_21\:DS_Offset = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_21\:Ref_Filename = "SM_OPER_AUX_OTT3F__20210624T082406_20500101T000000_700_001_1" ;
		string :VH\:SPH\:LODS\:Data_Set_21\:Num_DSR = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_21\:DSR_Size = "00000000" ;
		string :VH\:SPH\:LODS\:Data_Set_21\:Byte_Order = "0000" ;
		string :VH\:SPH\:LODS\:Data_Set_22\:DS_Name = "DGGRFI_FILE" ;
		string :VH\:SPH\:LODS\:Data_Set_22\:DS_Type = "R" ;
		string :VH\:SPH\:LODS\:Data_Set_22\:DS_Size = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_22\:DS_Offset = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_22\:Ref_Filename = "SM_OPER_AUX_DGGRFI_20210629T000711_20500101T000000_600_001_1" ;
		string :VH\:SPH\:LODS\:Data_Set_22\:Num_DSR = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_22\:DSR_Size = "00000000" ;
		string :VH\:SPH\:LODS\:Data_Set_22\:Byte_Order = "0000" ;
		string :VH\:SPH\:LODS\:Data_Set_23\:DS_Name = "MIXED_SCENE_OTT_FILE" ;
		string :VH\:SPH\:LODS\:Data_Set_23\:DS_Type = "R" ;
		string :VH\:SPH\:LODS\:Data_Set_23\:DS_Size = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_23\:DS_Offset = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_23\:Ref_Filename = "SM_OPER_AUX_MSOTT__20050101T000000_20500101T000000_001_002_3" ;
		string :VH\:SPH\:LODS\:Data_Set_23\:Num_DSR = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_23\:DSR_Size = "00000000" ;
		string :VH\:SPH\:LODS\:Data_Set_23\:Byte_Order = "0000" ;
		string :VH\:SPH\:L2PL\:Start_Lat = "-075.538036" ;
		string :VH\:SPH\:L2PL\:Start_Long = "-094.410663" ;
		string :VH\:SPH\:L2PL\:Stop_Lat = "+081.601490" ;
		string :VH\:SPH\:L2PL\:Stop_Long = "+017.400949" ;
		string :VH\:SPH\:L2PL\:Mid_Lat = "-005.823823" ;
		string :VH\:SPH\:L2PL\:Mid_Lon = "+114.700199" ;
		string :VH\:SPH\:L2PL\:Southernmost_Latitude = "-063.270000" ;
		string :VH\:SPH\:L2PL\:Southernmost_Gridpoint_ID = "7240286" ;
		string :VH\:SPH\:L2PL\:Northernmost_Latitude = "+080.555000" ;
		string :VH\:SPH\:L2PL\:Northernmost_Gridpoint_ID = "4094657" ;
		string :VH\:SPH\:L2PL\:Easternmost_Longitude = "+148.524002" ;
		string :VH\:SPH\:L2PL\:Easternmost_Gridpoint_ID = "7243351" ;
		string :VH\:SPH\:L2PL\:Westernmost_Longitude = "+023.934000" ;
		string :VH\:SPH\:L2PL\:Westernmost_Gridpoint_ID = "4081389" ;
		string :VH\:MPH\:Ref_Doc = "SO-TN-IDR-GS-0006" ;
		string :VH\:MPH\:Acquisition_Station = "SVLD" ;
		string :VH\:MPH\:Processing_Centre = "ESAC" ;
		string :VH\:MPH\:Logical_Proc_Centre = "FPC" ;
		string :VH\:MPH\:Product_Confidence = "NOMINAL" ;
		string :VH\:MPH\:OI\:Phase = "+001" ;
		string :VH\:MPH\:OI\:Cycle = "+037" ;
		string :VH\:MPH\:OI\:Rel_Orbit = "+01161" ;
		string :VH\:MPH\:OI\:Abs_Orbit = "+61281" ;
		string :VH\:MPH\:OI\:OSV_TAI = "TAI=2021-06-30T21:58:37.000000" ;
		string :VH\:MPH\:OI\:OSV_UTC = "UTC=2021-06-30T21:58:00.000000" ;
		string :VH\:MPH\:OI\:OSV_UT1 = "UT1=2021-06-30T21:58:00.590000" ;
		string :VH\:MPH\:OI\:X_Position = "+0146839.075" ;
		string :VH\:MPH\:OI\:Y_Position = "-2215887.397" ;
		string :VH\:MPH\:OI\:Z_Position = "-6791787.132" ;
		string :VH\:MPH\:OI\:X_Velocity = "-4093.431900" ;
		string :VH\:MPH\:OI\:Y_Velocity = "+5989.437140" ;
		string :VH\:MPH\:OI\:Z_Velocity = "-2043.308610" ;
		string :VH\:MPH\:OI\:Vector_Source = "FP" ;
		:history = "Mon Sep 25 18:37:41 2023: ncks -d n_grid_points,100,92700,1800 /scratch1/NCEPDEV/stmp4/Shastri.Paturi/forAndrew/gdas.20210701/00/SSS/SM_OPER_MIR_OSUDP2_20210630T215911_20210630T225230_700_001_1.nc sss_smos_2.nc" ;
		:NCO = "netCDF Operators version 5.0.6 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco)" ;
data:

 A_card = _, _, _, _, _, _, _, _, 47.73457, 49.38494, _, 51.50238, 48.75237, 
    49.85275, 50.02007, 52.50782, 50.81105, 48.75327, 54.03027, _, 53.25703, 
    _, _, _, 58.30848, 58.91204, 60.08769, 60.46875, _, _, _, 59.17318, 
    57.85364, _, _, _, _, _, _, 23.93925, _, _, _, _, _, _, 48.02232, 
    48.59546, 26.67431, _, 48.07984, _ ;

 Coast_distance = 4, 2, 20, _, 12, 15, 8, 16, 53, 62, 48, 39, 80, 55, 55, 57, 
    32, 44, 5, 28, 11, _, 1, _, 18, 24, 22, 6, _, 1, _, 2, 3, 1, _, 3, 5, _, 
    2, 3, _, 16, _, _, _, 1, 3, 10, 5, 4, 14, 30 ;

 Control_Flags_Acard = 51548168, 437420040, 453122049, 50468865, 437420040, 
    163840, 168984584, 16945152, 8814592, 8815104, 50468865, 59150344, 
    8815104, 59150864, 8815104, 8815104, 8815104, 8815104, 8815104, 
    453122049, 411468288, 50466817, 184680449, 50468865, 411468288, 
    411468288, 8815104, 25596416, 50462721, 50462721, 50468865, 8815104, 
    411468544, 50466817, 50468865, 453122048, 453122048, 50468865, 453122048, 
    446071560, 50468865, 453122049, 50468865, 50468865, 184680449, 453115905, 
    143032320, 411467776, 462852616, 34766856, 411467776, 453122049 ;

 Control_Flags_anom = 50499584, 520257536, 520230913, 50468865, 453148672, 
    50495488, 184713216, 50499584, 8814592, 8815104, 50468865, 59674650, 
    8815104, 59675184, 8815104, 8815104, 8815104, 8815136, 8815136, 
    520230913, 478577152, 117575681, 184680449, 50468865, 445022768, 
    411468288, 8815136, 26120736, 117571585, 50462721, 50468865, 8815104, 
    478577440, 50466817, 50468865, 520271872, 520271872, 50468865, 520271872, 
    528918334, 50468865, 520230913, 50468865, 50468865, 184680449, 453115905, 
    143032320, 445023232, 462344732, 50495488, 411467776, 453122049 ;

 Control_Flags_corr = 50499584, 520257536, 520230913, 50468865, 453148672, 
    50495488, 184713216, 50499584, 8814592, 8815104, 50468865, 59674650, 
    8815104, 59675184, 8815104, 8815104, 8815104, 8815136, 8815136, 
    520230913, 478577152, 117575681, 184680449, 50468865, 445022768, 
    411468288, 8815136, 26120736, 117571585, 50462721, 50468865, 8815104, 
    478577440, 50466817, 50468865, 520271872, 520271872, 50468865, 520271872, 
    528918334, 50468865, 520230913, 50468865, 50468865, 184680449, 453115905, 
    143032320, 445023232, 462344732, 50495488, 411467776, 453122049 ;

 Control_Flags_uncorr = 50466816, 520224768, 520230913, 50468865, 453115904, 
    50462720, 184680448, 50466816, 8814592, 8814592, 50468865, 59150362, 
    8814592, 59150384, 8814592, 8814592, 8814592, 8814624, 8814624, 
    520230913, 478576640, 117575681, 184680449, 50468865, 445022256, 
    411467776, 8814624, 25595936, 117571585, 50462721, 50468865, 8814592, 
    478576928, 50466817, 50468865, 520239104, 520239104, 50468865, 520239104, 
    528917820, 50468865, 520230913, 50468865, 50468865, 184680449, 453115905, 
    143032320, 445023232, 461819932, 50462720, 411467776, 453122049 ;

 Dg_RFI_L1 = 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 10, 17, 3, 0, 23, 36, 0, 15, 110, 5, 0, 191, 191, 0, 204, 219, 
    0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 Dg_RFI_X = 0, 61, 6, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 4, 0, 34, 1, 16, 
    12, 0, 0, 0, 0, 0, 0, 24, 29, 0, 7, 64, 5, 0, 117, 113, 0, 112, 101, 0, 
    3, 0, 0, 7, 7, 3, 4, 0, 0, 1, 0 ;

 Dg_RFI_Y = 0, 59, 6, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 2, 0, 32, 2, 13, 
    12, 0, 0, 0, 0, 0, 0, 24, 27, 0, 9, 61, 4, 0, 118, 111, 0, 111, 106, 0, 
    2, 0, 0, 8, 6, 3, 5, 0, 0, 2, 0 ;

 Dg_RFI_probability = 1, 2, 9, 0, 4, 2, 2, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 
    0, 2, 11, 0, 2, 0, 3, 3, 1, 0, 1, 1, 0, 1, 4, 2, 0, 10, 12, 0, 16, 20, 0, 
    81, 0, 0, 2, 2, 2, 28, 3, 2, 24, 77 ;

 Dg_Suspect_ice = _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, 140, _, _, 16, _, _, _ ;

 Dg_af_fov = _, 150, _, _, 145, 172, _, _, 150, 57, _, _, 168, _, 167, _, 
    157, _, 173, _, _, _, _, _, 147, 163, 1, _, 16, 159, _, 2, 148, _, _, 
    149, 165, _, 167, 150, _, _, _, _, 150, 29, 163, 162, _, _, _, _ ;

 Dg_border_fov = 11, 30, 9, _, 30, 26, 9, 8, 30, 28, 2, 8, 16, 10, 25, 13, 
    14, 9, 35, 5, 11, 9, 8, _, 32, 17, 13, 9, 60, 54, _, 13, 32, 11, _, 31, 
    17, _, 35, 27, _, 5, _, _, 32, 105, 14, 28, 10, 9, 10, 2 ;

 Dg_chi2_Acard = 174, 267, _, _, 563, 117, 230, 124, 113, 97, _, 147, 111, 
    51, 113, 114, 111, 101, 103, _, 89, _, _, _, 120, 88, 95, 83, _, _, _, 
    99, 103, _, _, _, _, _, _, 8780, _, _, _, _, _, _, 116, 112, 186, 179, 
    118, _ ;

 Dg_chi2_P_Acard = 993, 1000, _, _, 1000, 967, 1000, 845, 917, 386, _, 965, 
    894, 24, 906, 811, 877, 545, 621, _, 318, _, _, _, 976, 82, 382, 281, _, 
    _, _, 497, 589, _, _, _, _, _, _, 1000, _, _, _, _, _, _, 954, 908, 993, 
    999, 868, _ ;

 Dg_chi2_P_corr = _, _, _, _, _, _, _, _, 897, 322, _, 950, 882, 2, 867, 784, 
    859, 497, 571, _, 170, _, _, _, 971, 72, 310, 201, _, _, _, 456, 244, _, 
    _, _, _, _, _, 1000, _, _, _, _, _, _, 947, 823, 1000, _, 853, _ ;

 Dg_chi2_P_uncorr = _, _, _, _, _, _, _, _, 897, 327, _, 950, 891, 1, 830, 
    806, 933, 563, 892, _, 187, _, _, _, 998, 166, 448, 186, _, _, _, 821, 
    498, _, _, _, _, _, _, 1000, _, _, _, _, _, _, 947, 823, 1000, _, 853, _ ;

 Dg_chi2_corr = _, _, _, _, _, _, _, _, 112, 95, _, 142, 111, 37, 111, 112, 
    110, 98, 102, _, 80, _, _, _, 119, 87, 93, 77, _, _, _, 98, 90, _, _, _, 
    _, _, _, 9485, _, _, _, _, _, _, 115, 109, 1232, _, 116, _ ;

 Dg_chi2_uncorr = _, _, _, _, _, _, _, _, 112, 95, _, 142, 111, 37, 109, 113, 
    114, 102, 113, _, 81, _, _, _, 131, 91, 98, 76, _, _, _, 113, 99, _, _, 
    _, _, _, _, 11693, _, _, _, _, _, _, 115, 109, 5016, _, 116, _ ;

 Dg_galactic_Noise_Error = _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _ ;

 Dg_moonglint = _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _ ;

 Dg_num_iter_Acard = 4, 6, _, _, 7, 7, 5, 6, 7, 7, _, 6, 7, 6, 7, 6, 7, 6, 7, 
    _, 6, _, _, _, 7, 7, 7, 6, _, _, _, 6, 7, _, _, _, _, _, _, 5, _, _, _, 
    _, _, _, 7, 7, 6, 4, 6, _ ;

 Dg_num_iter_corr = _, _, _, _, _, _, _, _, 3, 2, _, 2, 2, 3, 3, 3, 3, 2, 3, 
    _, 3, _, _, _, 9, 2, 2, 2, _, _, _, 2, 6, _, _, _, _, _, _, 20, _, _, _, 
    _, _, _, 11, 20, 17, _, 2, _ ;

 Dg_num_iter_uncorr = _, _, _, _, _, _, _, _, 3, 2, _, 2, 2, 3, 3, 3, 3, 2, 
    2, _, 2, _, _, _, 3, 2, 2, 2, _, _, _, 3, 5, _, _, _, _, _, _, 20, _, _, 
    _, _, _, _, 11, 20, 7, _, 2, _ ;

 Dg_num_meas_l1c = 35, 235, 12, _, 233, 238, 63, 34, 240, 234, 2, 34, 228, 
    28, 228, 74, 219, 40, 231, 5, 69, 53, 43, _, 233, 223, 90, 30, 138, 218, 
    _, 88, 240, 30, _, 235, 224, _, 223, 237, _, 5, _, _, 240, 210, 223, 233, 
    28, 43, 75, 2 ;

 Dg_num_meas_valid = 24, 66, _, _, 158, 185, 54, 26, 170, 154, _, 26, 192, 
    18, 170, 61, 180, 31, 131, _, 34, 26, 35, _, 163, 191, 77, 21, 49, 103, 
    _, 69, 75, 16, _, _, _, _, _, 32, _, _, _, _, 159, 90, 188, 176, 18, 34, 
    62, _ ;

 Dg_quality_SSS_anom = 0, 0, 0, 0, 0, 0, 0, 0, 247, 300, 0, 0, 125, _, 131, 
    298, 92, 306, 116, 0, 219, 0, 0, 0, _, 57, 154, 210, 0, 0, 0, 168, 128, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 288, _, _, 0, 472, 0 ;

 Dg_quality_SSS_corr = _, _, _, _, _, _, _, _, 247, 300, _, _, 125, _, 131, 
    298, 92, 306, 116, _, 219, _, _, _, _, 57, 154, 210, _, _, _, 168, 128, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, 288, _, _, _, 472, _ ;

 Dg_quality_SSS_uncorr = _, _, _, _, _, _, _, _, 247, 300, _, _, 125, _, 131, 
    298, 92, 306, 116, _, 219, _, _, _, _, 57, 154, 210, _, _, _, 168, 128, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, 288, _, _, _, 472, _ ;

 Dg_sky = 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 46, 0, 0, 0, 33, 0, 0, 33, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0 ;

 Dg_sun_glint_L2 = _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _ ;

 Dg_sun_glint_area = _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 5, _, 
    _, 83, _, _, _, _, 43, _, 2 ;

 Dg_sun_glint_fov = _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _ ;

 Dg_sun_tails = _, 59, _, _, 52, 16, 12, 9, 19, _, _, _, 16, 15, 192, 16, 19, 
    16, 15, 5, _, _, 1, _, 13, 25, 15, 6, 15, 17, _, 16, 86, 15, _, 15, 53, 
    _, 27, 99, _, _, _, _, 17, 15, 32, 158, 20, _, 17, _ ;

 Equiv_ftprt_diam = 56.89935, 56.06676, 63.05637, _, 57.97224, 51.55901, 
    50.19272, 56.48489, 55.55499, 60.5041, 66.63572, 56.59513, 48.7635, 
    57.84214, 51.72989, 48.60321, 48.40091, 51.88385, 50.17692, 64.95056, 
    48.58825, 51.28894, 53.06034, _, 54.72203, 47.95681, 46.54311, 55.8958, 
    57.44204, 48.42532, _, 46.30187, 52.61933, 55.7595, _, 53.0805, 48.17634, 
    _, 48.29556, 52.00186, _, 63.55217, _, _, 54.16161, 60.73178, 48.21849, 
    50.94963, 56.86495, 52.96722, 47.61303, 65.34607 ;

 Grid_Point_ID = 6251019, 7186392, 7194052, 7213054, 7233627, 7235697, 
    7235661, 7242327, 7258289, 7248082, 7261320, 7230646, 8109073, 8141853, 
    8094752, 8124977, 8090169, 8120903, 8087128, 8120929, 8066611, 8057411, 
    8052315, 8051827, 8072921, 8061140, 8046761, 8086249, 8068893, 8059160, 
    8042776, 8040189, 8039228, 8030983, 8071506, 8049538, 8035708, 8027528, 
    8037286, 8022951, 8041944, 8059331, 4045749, 4065379, 4084876, 4066467, 
    4080816, 4078787, 4055194, 4102838, 4072659, 4120306 ;

 Latitude = -76.151, -77.41, -74.643, -71.861, -64.609, -63.034, -64.906, 
    -63.205, -55.638, -54.537, -57.479, -58.616, -48.685, -51.452, -44.391, 
    -46.513, -40.182, -42.866, -35.332, -39.175, -37.132, -33.301, -28.93, 
    -25.44, -14.805, -13.467, -16.861, -14.725, -4.935, -4.42, -2.378, 
    -5.508, 2.697, -3.076, 1.48, 10.232, 11.234, 13.737, 16.148, 18.106, 
    22.444, 17.864, 51.638, 69.291, 74.944, 74.356, 77.42, 77.959, 71.973, 
    80.454, 76.93, 87.38 ;

 Longitude = -157.126, 177.916, -170.177, 165.449, 143.108, 138.427, 147.869, 
    148.091, 134.345, 123.998, 144.011, 120.997, 126.188, 137.108, 122.752, 
    131.805, 122.686, 131.029, 123.431, 131.595, 117.177, 115.688, 114.405, 
    114.364, 119.251, 116.545, 113.311, 122.324, 117.944, 115.496, 111.48, 
    110.942, 110.625, 108.663, 118.323, 113.515, 110.075, 108.134, 110.859, 
    107.175, 112.003, 116.105, 101.016, 82.105, 85.012, 60.59, 64.585, 
    51.372, 58.422, 86.772, 37.611, 56.383 ;

 Mean_acq_time = 7851.918, 7851.919, 7851.919, _, 7851.922, 7851.922, 
    7851.922, 7851.922, 7851.924, 7851.924, 7851.923, 7851.924, 7851.925, 
    7851.925, 7851.926, 7851.926, 7851.927, 7851.927, 7851.928, 7851.927, 
    7851.928, 7851.929, 7851.93, _, 7851.932, 7851.932, 7851.932, 7851.932, 
    7851.934, 7851.934, _, 7851.935, 7851.936, 7851.935, _, 7851.937, 
    7851.937, _, 7851.938, 7851.938, _, 7851.938, _, _, 7851.95, 7851.95, 
    7851.951, 7851.951, 7851.951, 7851.951, 7851.952, 7851.952 ;

 SSS_anom = _, _, _, _, _, _, _, _, 1.628859, 1.243454, _, _, -4.30769, _, 
    -2.113121, _, -4.591354, _, -0.1896324, _, _, _, _, _, -1.178625, 
    -1.055939, 0.1436996, _, _, _, _, -0.2785378, 0.04353333, _, _, _, _, _, 
    _, -30.69485, _, _, _, _, _, _, 0.1373024, 2.33411, _, _, _, _ ;

 SSS_climatology = 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 
    2897, 3320, 65535, 65535, 3392, 65535, 3489, 65535, 3511, 65535, 3614, 
    65535, 65535, 65535, 65535, 65535, 3216, 3425, 3540, 65535, 65535, 65535, 
    65535, 3238, 2912, 65535, 65535, 65535, 65535, 65535, 65535, 3328, 65535, 
    65535, 65535, 65535, 65535, 65535, 3139, 2889, 65535, 65535, 65535, 65535 ;

 SSS_corr = _, _, _, _, _, _, _, _, 30.59692, 34.46416, _, _, 29.57378, 
    33.6181, 32.66331, 38.32122, 30.43209, 28.0537, 35.61701, _, 33.53222, _, 
    _, _, 32.95224, 33.26748, 34.88172, 34.5612, _, _, _, 32.28378, 31.75333, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, 31.5253, 31.22411, 0.9942121, _, 
    33.04895, _ ;

 SSS_uncorr = _, _, _, _, _, _, _, _, 30.59486, 34.44645, _, _, 29.61531, 
    33.32262, 32.77388, 38.15655, 30.52065, 26.85291, 35.95137, _, 33.39886, 
    _, _, _, 30.98137, 33.19106, 35.5447, 33.2958, _, _, _, 32.10446, 
    29.16653, _, _, _, _, _, _, 2.586151, _, _, _, _, _, _, 31.5253, 
    31.22411, 0.9942121, _, 33.04895, _ ;

 SST = _, _, _, _, _, _, _, _, 2.82431, 3.93631, _, 1.423431, 7.957458, 
    5.960266, 9.887207, 9.335083, 12.49179, 11.07925, 15.82275, _, 17.14066, 
    _, _, _, 27.30756, 27.66653, 26.68677, 27.69809, _, _, _, 29.53842, 
    29.60687, _, _, _, _, _, _, 29.82776, _, _, _, _, _, _, 0.6308899, 
    0.7425537, 0.4602051, _, 0.1035767, _ ;

 Science_Flags_Acard = 2109467, 2234779, 14745, 4208640, 2111897, 70041, 
    2111899, 12441, 20737, 12673, 70017, 12673, 39041, 39041, 15489, 39041, 
    15489, 15489, 15747, 40065, 23937, 4217858, 73474, 4209920, 72449, 72577, 
    72449, 72451, 37762, 37634, 4208128, 70403, 20995, 13058, 4217344, 37635, 
    37763, 4208384, 13187, 136067, 4209408, 37761, 4202496, 4203520, 8218, 
    16426, 20491, 69641, 69675, 2105627, 135561, 12569 ;

 Science_Flags_anom = 12315, 137627, 14745, 4208640, 14745, 70041, 14747, 
    12441, 20737, 12673, 70017, 12673, 39041, 39041, 15489, 39041, 15489, 
    15489, 15747, 40065, 23937, 4217858, 73474, 4209920, 72449, 72577, 72449, 
    72451, 37762, 37634, 4208128, 70403, 20995, 13058, 4217344, 37635, 37763, 
    4208384, 13187, 136067, 4209408, 37761, 4202496, 4203520, 8218, 16426, 
    20491, 69641, 69675, 8475, 135561, 12569 ;

 Science_Flags_corr = 12315, 137627, 14745, 4208640, 14745, 70041, 14747, 
    12441, 20737, 12673, 70017, 12673, 39041, 39041, 15489, 39041, 15489, 
    15489, 15747, 40065, 23937, 4217858, 73474, 4209920, 72449, 72577, 72449, 
    72451, 37762, 37634, 4208128, 70403, 20995, 13058, 4217344, 37635, 37763, 
    4208384, 13187, 136067, 4209408, 37761, 4202496, 4203520, 8218, 16426, 
    20491, 69641, 69675, 8475, 135561, 12569 ;

 Science_Flags_uncorr = 12315, 137627, 14745, 4208640, 14745, 70041, 14747, 
    12441, 20737, 12673, 70017, 12673, 39041, 39041, 15489, 39041, 15489, 
    15489, 15747, 40065, 23937, 4217858, 73474, 4209920, 72449, 72577, 72449, 
    72451, 37762, 37634, 4208128, 70403, 20995, 13058, 4217344, 37635, 37763, 
    4208384, 13187, 136067, 4209408, 37761, 4202496, 4203520, 8218, 16426, 
    20491, 69641, 69675, 8475, 135561, 12569 ;

 Sigma_Acard = _, _, _, _, _, _, _, _, 0.5851961, 0.5876574, _, 1.735356, 
    0.5692883, 1.606627, 0.6001664, 0.9319488, 0.5823345, 1.144666, 
    0.6193509, _, 1.104503, _, _, _, 0.7022212, 0.5980276, 0.8724535, 
    1.986215, _, _, _, 0.9349416, 0.7858232, _, _, _, _, _, _, 6.679135, _, 
    _, _, _, _, _, 0.5980026, 0.6083651, 1.178608, _, 0.9472713, _ ;

 Sigma_SSS_anom = _, _, _, _, _, _, _, _, 1.943289, 2.015971, _, _, 2.21241, 
    4.420088, 2.091019, 3.159312, 1.382608, 2.935465, 1.132476, _, 1.895663, 
    _, _, _, 0.6969603, 0.5503999, 0.8192711, 1.835188, _, _, _, 0.8325468, 
    0.6733742, _, _, _, _, _, _, _, _, _, _, _, _, _, 2.208032, 2.230621, 
    213.0026, _, 3.79549, _ ;

 Sigma_SSS_corr = _, _, _, _, _, _, _, _, 1.943289, 2.015971, _, _, 2.21241, 
    4.420088, 2.091019, 3.159312, 1.382608, 2.935465, 1.132476, _, 1.895663, 
    _, _, _, 0.6969603, 0.5503999, 0.8192711, 1.835188, _, _, _, 0.8325468, 
    0.6733742, _, _, _, _, _, _, _, _, _, _, _, _, _, 2.208032, 2.230621, 
    213.0026, _, 3.79549, _ ;

 Sigma_SSS_uncorr = _, _, _, _, _, _, _, _, 1.943316, 2.016585, _, _, 
    2.214404, 4.432564, 2.068832, 3.181352, 1.313231, 3.020818, 1.194507, _, 
    1.831774, _, _, _, 0.6450708, 0.4912785, 0.8267764, 1.813485, _, _, _, 
    0.8847318, 0.6245384, _, _, _, _, _, _, 90.83298, _, _, _, _, _, _, 
    2.208032, 2.230621, 430.4953, _, 3.79549, _ ;

 Sigma_Tb_42_5H = _, _, _, _, _, _, _, _, 0.5803481, 0.7497043, _, _, 
    0.8924729, _, 1.074311, 1.408248, 0.7830504, 1.170192, 0.7262191, _, 
    1.017727, _, _, _, 0.6223353, 0.5363076, 0.6052372, _, _, _, _, 
    0.6366693, 0.6210805, _, _, _, _, _, _, 13.20704, _, _, _, _, _, _, 
    0.6847072, 0.9120925, _, _, 0.8533247, _ ;

 Sigma_Tb_42_5V = _, _, _, _, _, _, _, _, 0.6388904, 0.7884085, _, _, 
    1.023682, _, 1.144722, 1.602629, 0.8156266, 1.406483, 0.7618073, _, 
    1.191876, _, _, _, 0.6186877, 0.5079992, 0.6453832, _, _, _, _, 
    0.7107596, 0.6153561, _, _, _, _, _, _, 18.28141, _, _, _, _, _, _, 
    0.6457273, 0.7188643, _, _, 1.006405, _ ;

 Sigma_Tb_42_5X = _, _, _, _, _, _, _, _, 0.6142722, 0.7770153, _, _, 
    0.88337, _, 1.072063, 1.601871, 0.777356, 1.609143, 0.7344985, _, 
    1.363688, _, _, _, 0.8075515, 0.5317979, 0.9279311, _, _, _, _, 1.040271, 
    0.6366233, _, _, _, _, _, _, 13.61083, _, _, _, _, _, _, 0.6773354, 
    0.9011479, _, _, 1.110289, _ ;

 Sigma_Tb_42_5Y = _, _, _, _, _, _, _, _, 0.6539022, 0.7980523, _, _, 
    1.014643, _, 1.137706, 1.635368, 0.8100698, 1.565964, 0.7656733, _, 
    1.393147, _, _, _, 0.8108457, 0.5046097, 0.9314546, _, _, _, _, 1.05729, 
    0.63436, _, _, _, _, _, _, 17.56855, _, _, _, _, _, _, 0.6403679, 
    0.7292545, _, _, 1.134751, _ ;

 Sigma_WS_corr = _, _, _, _, _, 2803, 2577, 2512, 2597, 2627, 2515, 2817, 
    2367, 2819, 2426, 2784, 2510, 2814, 2509, 2816, 2815, 2822, 2806, 2763, 
    2608, 2511, 2800, 2813, 2592, 2594, 2822, 2809, 2642, 2805, 2819, 2821, 
    2821, 2821, 2821, 2817, 2828, 2828, 2721, 2721, 2721, 2520, 2226, 2226, 
    2811, 2760, 2811, 2823 ;

 Tb_42_5H = _, _, _, _, _, _, _, _, 78.74249, 79.03468, _, _, 83.72257, _, 
    82.71999, 80.91987, 81.44019, 82.46483, 79.64092, _, 80.06966, _, _, _, 
    78.75982, 78.64634, 77.13834, _, _, _, _, 78.37289, 79.25348, _, _, _, _, 
    _, _, 96.80058, _, _, _, _, _, _, 76.31535, 75.99258, _, _, 78.17581, _ ;

 Tb_42_5V = _, _, _, _, _, _, _, _, 121.9867, 121.698, _, _, 126.7233, _, 
    125.5164, 123.1936, 125.1497, 126.2615, 122.7925, _, 123.7155, _, _, _, 
    123.227, 123.0001, 121.4938, _, _, _, _, 123.3869, 124.1231, _, _, _, _, 
    _, _, 147.2917, _, _, _, _, _, _, 120.3693, 120.3368, _, _, 120.8457, _ ;

 Tb_42_5X = _, _, _, _, _, _, _, _, 86.6127, 89.21529, _, _, 85.59736, _, 
    86.38583, 100.1518, 83.64706, 110.5141, 82.85757, _, 99.1396, _, _, _, 
    86.37729, 80.57986, 94.36686, _, _, _, _, 94.69478, 86.5731, _, _, _, _, 
    _, _, 103.6411, _, _, _, _, _, _, 78.37074, 80.48462, _, _, 96.19685, _ ;

 Tb_42_5Y = _, _, _, _, _, _, _, _, 117.4025, 114.8389, _, _, 128.0181, _, 
    125.1165, 107.1409, 126.2634, 101.4164, 122.9822, _, 108.045, _, _, _, 
    119.0049, 124.4646, 107.7274, _, _, _, _, 110.4799, 120.208, _, _, _, _, 
    _, _, 143.4219, _, _, _, _, _, _, 121.7208, 119.2336, _, _, 106.1588, _ ;

 WS = _, _, _, _, _, _, _, _, 6.862242, 11.02606, _, 10.45476, 18.95231, 
    13.11163, 17.19608, 16.74842, 14.2471, 14.34991, 11.38515, _, 10.94148, 
    _, _, _, 6.50735, 7.431638, 4.760453, 3.806333, _, _, _, 4.937733, 
    2.75331, _, _, _, _, _, _, 8.910588, _, _, _, _, _, _, 1.762767, 
    2.880984, 2.587532, _, 9.089414, _ ;

 WS_corr = _, _, _, _, _, 11210, 8480, 4481, 7436, 11017, 11057, 8794, 18619, 
    12899, 17727, 17515, 12660, 13852, 12381, 12708, 11290, 9616, 6069, 6028, 
    7241, 7723, 4781, 3768, 8134, 7634, 8733, 4680, 6159, 4186, 4655, 4446, 
    4446, 4446, 4446, 20535, 37953, 32911, 21054, 21054, 21054, 2434, 925, 
    129, 6223, 329, 8763, 9906 ;

 X_swath = -597.8799, -266.4582, _, _, -303.0927, -171.526, -483.2304, 
    -593.0931, -268.8257, 328.2765, _, 596.4514, 24.21224, -613.5121, 
    163.3268, -450.7834, 60.41842, -525.3317, -133.4874, _, 458.3513, _, _, 
    _, -267.2321, -15.27115, 402.6631, -591.2664, _, _, _, 399.5669, 
    241.3157, _, _, -248.7068, 95.24609, _, -104.8272, 229.7502, _, _, _, _, 
    _, _, 32.41647, 184.4597, 603.1434, -545.4169, 434.0908, _ ;
}
