netcdf rads_adt_c2_2018105.tmp {
dimensions:
	time = UNLIMITED ; // (11 currently)
variables:
	int adt_egm2008(time) ;
		adt_egm2008:_FillValue = 2147483647 ;
		adt_egm2008:long_name = "absolute dynamic topography (EGM2008)" ;
		adt_egm2008:standard_name = "absolute_dynamic_topography_egm2008" ;
		adt_egm2008:units = "m" ;
		adt_egm2008:scale_factor = 0.0001 ;
		adt_egm2008:coordinates = "lon lat" ;
	int adt_xgm2016(time) ;
		adt_xgm2016:_FillValue = 2147483647 ;
		adt_xgm2016:long_name = "absolute dynamic topography (XGM2016)" ;
		adt_xgm2016:standard_name = "absolute_dynamic_topography_xgm2016" ;
		adt_xgm2016:units = "m" ;
		adt_xgm2016:scale_factor = 0.0001 ;
		adt_xgm2016:coordinates = "lon lat" ;
	int cycle(time) ;
		cycle:_FillValue = 2147483647 ;
		cycle:long_name = "cycle number" ;
		cycle:field = 9905s ;
	int lat(time) ;
		lat:_FillValue = 2147483647 ;
		lat:long_name = "latitude" ;
		lat:standard_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:scale_factor = 1.e-07 ;
		lat:field = 201s ;
		lat:comment = "Positive latitude is North latitude, negative latitude is South latitude" ;
	int lon(time) ;
		lon:_FillValue = 2147483647 ;
		lon:long_name = "longitude" ;
		lon:standard_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:scale_factor = 1.e-07 ;
		lon:field = 301s ;
		lon:comment = "East longitude relative to Greenwich meridian" ;
	int pass(time) ;
		pass:_FillValue = 2147483647 ;
		pass:long_name = "pass number" ;
		pass:field = 9906s ;
	short sla(time) ;
		sla:_FillValue = 32767s ;
		sla:long_name = "sea level anomaly" ;
		sla:standard_name = "sea_surface_height_above_sea_level" ;
		sla:units = "m" ;
		sla:quality_flag = "swh sig0 range_rms range_numval flags peakiness" ;
		sla:scale_factor = 0.0001 ;
		sla:coordinates = "lon lat" ;
		sla:field = 0s ;
		sla:comment = "Sea level determined from satellite altitude - range - all altimetric corrections" ;
	double time_mjd(time) ;
		time_mjd:long_name = "Modified Julian Days" ;
		time_mjd:standard_name = "time" ;
		time_mjd:units = "days since 1858-11-17 00:00:00 UTC" ;
		time_mjd:field = 105s ;
		time_mjd:comment = "UTC time of measurement expressed in Modified Julian Days" ;

// global attributes:
		:Conventions = "CF-1.7" ;
		:title = "RADS 4 pass file" ;
		:institution = "EUMETSAT / NOAA / TU Delft" ;
		:source = "radar altimeter" ;
		:references = "RADS Data Manual, Version 4.2 or later" ;
		:featureType = "trajectory" ;
		:ellipsoid = "TOPEX" ;
		:ellipsoid_axis = 6378136.3 ;
		:ellipsoid_flattening = 0.00335281317789691 ;
		:filename = "rads_adt_c2_2018105.nc" ;
		:mission_name = "CRYOSAT2" ;
		:mission_phase = "a" ;
		:log01 = "2019-01-11 | rads2nc --ymd=180415000000,180416000000 -C1,1000 -Sc2 -Vadt_egm2008,adt_xgm2016,sla,time_mjd,lon,lat,cycle,pass -Xxgm2016 -Xadt.xml -o/ftp/rads/adt//2018/rads_adt_c2_2018105.nc: RAW data from" ;
		:history = "Fri Jan 26 15:41:52 2024: ncks -d time,0,10 /scratch1/NCEPDEV/stmp4/Shastri.Paturi/forAndrew/gdas.20180415/00/adt/rads_adt_c2_2018105.nc rads_adt_c2_2018105.tmp.nc\n",
			"2019-01-11 12:29:43 : rads2nc --ymd=180415000000,180416000000 -C1,1000 -Sc2 -Vadt_egm2008,adt_xgm2016,sla,time_mjd,lon,lat,cycle,pass -Xxgm2016 -Xadt.xml -o/ftp/rads/adt//2018/rads_adt_c2_2018105.nc" ;
		:NCO = "netCDF Operators version 5.0.6 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco)" ;
data:

 adt_egm2008 = 6867, 6893, 6974, 6663, 6528, 6809, 7148, 6855, 6633, 6939, 
    7166 ;

 adt_xgm2016 = 5783, 6037, 6465, 6345, 6508, 6956, 7245, 6694, 6292, 6668, 
    6589 ;

 cycle = 104, 104, 104, 104, 104, 104, 104, 104, 104, 104, 104 ;

 lat = 202161175, 201588349, 201015521, 200442691, 199869857, 199297020, 
    198724180, 198151338, 197578493, 197005645, 196432796 ;

 lon = -1070968218, -1071030446, -1071092657, -1071154851, -1071217028, 
    -1071279190, -1071341335, -1071403463, -1071465575, -1071527671, 
    -1071589751 ;

 pass = 314, 314, 314, 314, 314, 314, 314, 314, 314, 314, 314 ;

 sla = -699, -484, -401, -699, -937, -621, -503, -456, -738, -583, -148 ;

 time_mjd = 58223.0000057087, 58223.0000166281, 58223.0000275475, 
    58223.0000384669, 58223.0000493863, 58223.0000603057, 58223.0000712251, 
    58223.0000821446, 58223.000093064, 58223.0001039834, 58223.0001149028 ;
}
