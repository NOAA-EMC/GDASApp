netcdf viirs_aod {
dimensions:
	Rows = 10 ;
	Columns = 10 ;
variables:
	float AOD550(Rows, Columns) ;
		AOD550:long_name = "Aerosol optical depth at 550 nm" ;
		AOD550:coordinates = "Longitude Latitude" ;
		AOD550:units = "1" ;
		AOD550:_FillValue = -999.999f ;
		AOD550:valid_range = -0.05f, 5.f ;
	float Latitude(Rows, Columns) ;
		Latitude:long_name = "Latitude" ;
		Latitude:units = "degrees_north" ;
		Latitude:comments = "Pixel latitude in field Latitude (degree)" ;
		Latitude:_FillValue = -999.f ;
		Latitude:valid_range = -90.f, 90.f ;
	float Longitude(Rows, Columns) ;
		Longitude:long_name = "Longitude" ;
		Longitude:units = "degrees_east" ;
		Longitude:comments = "Pixel longitude in field Longitude (degree)" ;
		Longitude:_FillValue = -999.f ;
		Longitude:valid_range = -180.f, 180.f ;
	byte QCAll(Rows, Columns) ;
		QCAll:long_name = "Retrieval quality:  0: high; 1: medium; 2: low; 3: no retrieval" ;
		QCAll:coordinates = "Longitude Latitude" ;
		QCAll:units = "1" ;
		QCAll:_FillValue = -128b ;
		QCAll:valid_range = 0b, 3b ;
	byte QCPath(Rows, Columns) ;
		QCPath:long_name = "Flags for retrieval path (0-No/1-Yes): bit 0: retrieval over water; bit 1: over bright land; bit 2: over glint water; bit 3: retrieval with SW scheme over land; bit 4: retrieval with SWIR scheme over land; bit 5: retrieval over bright-land algorithm" ;
		QCPath:coordinates = "Longitude Latitude" ;
		QCPath:units = "1" ;
		QCPath:_FillValue = -128b ;
		QCPath:valid_range = 0b, 31b ;
	float Residual(Rows, Columns) ;
		Residual:long_name = "Retrieval residual of the best solution" ;
		Residual:coordinates = "Longitude Latitude" ;
		Residual:units = "1" ;
		Residual:_FillValue = -999.999f ;
		Residual:valid_range = 0.f, 999.f ;

// global attributes:
		:Conventions = "CF-1.5" ;
		:Metadata_Conventions = "CF-1.5, Unidata Dataset Discovery v1.0" ;
		:standard_name_vocabulary = "CF Standard Name Table (version 17, 24 March 2011)" ;
		:project = "S-NPP Data Exploitation" ;
		:institution = "DOC/NOAA/NESDIS/NDE->S-NPP Data Exploitation, NESDIS, NOAA, U.S. Department of Commerce" ;
		:naming_authority = "gov.noaa.nesdis.nde" ;
		:satellite_name = "NPP" ;
		:instrument_name = "VIIRS" ;
		:title = "JPSS Risk Reduction Unique Aerosol Optical Depth" ;
		:summary = "Aerosol Optical Depth" ;
		:history = "Tue May 19 10:48:26 2020: ncks -v Latitude,Longitude,AOD550,QCPath,Residual,QCAll -d Columns,337,346 -d Rows,268,277 sample_viirs_class.nc sample_subset_testcase.nc\nVIIRS AOD Version 1.0" ;
		:processing_level = "NOAA Level 2" ;
		:references = "" ;
		:id = "ad1a951f-cc67-45d5-ab9d-b7be77d6a055" ;
		:Metadata_Link = "JRR-AOD_v1r1_npp_s201804150418347_e201804150419589_c201804150512090.nc" ;
		:start_orbit_number = 33494 ;
		:end_orbit_number = 33494 ;
		:day_night_data_flag = "day" ;
		:ascend_descend_data_flag = 0 ;
		:time_coverage_start = "2018-04-15T04:18:34Z" ;
		:time_coverage_end = "2018-04-15T04:19:58Z" ;
		:date_created = "2018-04-15T05:12:12Z" ;
		:cdm_data_type = "swath" ;
		:geospatial_first_scanline_first_fov_lat = 48.43998f ;
		:geospatial_first_scanline_last_fov_lat = 42.56979f ;
		:geospatial_last_scanline_first_fov_lat = 53.45447f ;
		:geospatial_last_scanline_last_fov_lat = 47.02182f ;
		:geospatial_first_scanline_first_fov_lon = 147.643f ;
		:geospatial_first_scanline_last_fov_lon = 108.7127f ;
		:geospatial_last_scanline_first_fov_lon = 147.7868f ;
		:geospatial_last_scanline_last_fov_lon = 105.0699f ;
		:geospatial_lat_units = "degrees_north" ;
		:geospatial_lon_units = "degrees_east" ;
		:geospatial_bounds = "POLYGON((147.643 48.44,108.713 42.5698,105.07 47.0218,147.787 53.4545,147.643 48.44))" ;
		:NCO = "netCDF Operators version 4.9.1 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco)" ;
data:

 AOD550 =
  0.08672047, 0.1280901, 0.01021459, 0.06967962, 0.1172924, 0.1077904, 
    0.0879033, 0.005564162, 0.05259846, 0.0844786,
  0.04495948, 0.07685012, 0.10102, 0.02387906, 0.007571651, 0.05067238, 
    0.01620957, 0.02683542, 0.1328741, 0.05480475,
  0.0328154, 0.1128744, 0.01603194, 0.1116905, 0.07046779, 0.08973835, 
    0.02214303, 0.02760522, 0.09676082, 0.007294201,
  0.03729188, 0.08136128, 0.034016, 0.05721173, 0.1383349, 0.1388035, 
    0.08501249, 0.08002064, 0.002229004, 0.1466849,
  0.08595434, 0.1187636, 0.0842336, 0.1316003, 0.08762938, 0.1063275, 
    0.02228002, 0.06426761, 0.1040835, 0.01569296,
  0.06594078, 0.02493032, 0.07604679, 0.1228554, 0.01351601, 0.1200103, 
    0.08476895, 0.08840216, 0.0297151, 0.06541774,
  0.04438556, 0.005633651, 0.004602726, 0.06796575, 0.1117296, 0.08359431, 
    0.05776704, 0.02521092, 0.1257392, 0.08985777,
  0.1174072, 0.1272764, 0.09047445, 0.1171591, 0.09236053, 0.003174779, 
    0.1125697, 0.02640632, 0.06877713, 0.07696841,
  0.07260314, 0.1266579, 0.02622208, 0.002195231, 0.1273146, 0.1114012, 
    0.06850463, 0.06253476, 0.01750943, 0.05080187,
  0.01419886, 0.1073746, 0.01156281, 0.03089254, 0.08606643, 0.04407473, 
    0.09835901, 0.1205353, 0.05268203, 0.01401606 ;

 Latitude =
  51.28726, 51.28702, 51.28678, 51.28655, 51.28631, 51.28606, 51.28583, 
    51.28558, 51.28534, 51.2851,
  51.299, 51.29874, 51.29851, 51.29826, 51.29802, 51.29776, 51.29752, 
    51.29727, 51.29702, 51.29676,
  51.31073, 51.31047, 51.31023, 51.30998, 51.30972, 51.30947, 51.30921, 
    51.30896, 51.3087, 51.30844,
  51.32247, 51.32221, 51.32196, 51.3217, 51.32143, 51.32117, 51.32091, 
    51.32065, 51.32038, 51.32011,
  51.25031, 51.25015, 51.24999, 51.24984, 51.24968, 51.24952, 51.24934, 
    51.24919, 51.24903, 51.24885,
  51.26204, 51.26187, 51.26171, 51.26155, 51.26138, 51.26121, 51.26104, 
    51.26087, 51.26069, 51.26053,
  51.27377, 51.27361, 51.27343, 51.27325, 51.27308, 51.27291, 51.27274, 
    51.27255, 51.27237, 51.27219,
  51.2855, 51.28532, 51.28515, 51.28497, 51.28478, 51.28461, 51.28442, 
    51.28424, 51.28405, 51.28386,
  51.29723, 51.29705, 51.29686, 51.29668, 51.29649, 51.2963, 51.29611, 
    51.29593, 51.29573, 51.29554,
  51.30896, 51.30877, 51.30858, 51.30839, 51.3082, 51.308, 51.3078, 51.30761, 
    51.30741, 51.30721 ;

 Longitude =
  142.8715, 142.8586, 142.8457, 142.8328, 142.82, 142.8071, 142.7943, 
    142.7815, 142.7687, 142.7559,
  142.8712, 142.8583, 142.8454, 142.8325, 142.8196, 142.8068, 142.794, 
    142.7811, 142.7684, 142.7556,
  142.8709, 142.858, 142.8451, 142.8322, 142.8193, 142.8065, 142.7937, 
    142.7808, 142.7681, 142.7553,
  142.8706, 142.8577, 142.8448, 142.8319, 142.819, 142.8062, 142.7933, 
    142.7805, 142.7677, 142.7549,
  142.8644, 142.8515, 142.8386, 142.8257, 142.8129, 142.8, 142.7872, 
    142.7744, 142.7617, 142.7489,
  142.864, 142.8511, 142.8382, 142.8253, 142.8125, 142.7997, 142.7868, 
    142.774, 142.7612, 142.7485,
  142.8637, 142.8508, 142.8379, 142.825, 142.8121, 142.7993, 142.7865, 
    142.7736, 142.7608, 142.7481,
  142.8633, 142.8504, 142.8375, 142.8246, 142.8118, 142.7989, 142.7861, 
    142.7733, 142.7605, 142.7477,
  142.8629, 142.85, 142.8371, 142.8242, 142.8114, 142.7985, 142.7857, 
    142.7729, 142.7601, 142.7473,
  142.8626, 142.8497, 142.8368, 142.8239, 142.811, 142.7981, 142.7853, 
    142.7725, 142.7597, 142.7469 ;

 QCAll =
  1, 0, 0, 0, 1, 2, 2, 2, 1, 2,
  2, 1, 2, 0, 1, 0, 1, 2, 1, 2,
  0, 2, 2, 2, 0, 2, 0, 1, 0, 0,
  1, 1, 2, 1, 2, 1, 0, 0, 1, 2,
  2, 0, 1, 1, 0, 1, 2, 1, 0, 2,
  1, 0, 1, 2, 1, 0, 0, 1, 0, 1,
  2, 0, 1, 0, 1, 0, 2, 2, 1, 2,
  0, 0, 1, 1, 2, 1, 1, 2, 0, 0,
  2, 2, 1, 2, 1, 0, 1, 1, 2, 1,
  2, 0, 0, 2, 1, 1, 2, 2, 2, 1 ;

 QCPath =
  1, 0, 1, 0, 1, 1, 1, 0, 1, 0,
  0, 0, 1, 0, 0, 0, 0, 0, 0, 1,
  1, 0, 0, 0, 1, 0, 1, 1, 1, 0,
  1, 0, 1, 1, 0, 0, 0, 1, 0, 0,
  1, 0, 0, 0, 0, 1, 0, 0, 1, 1,
  1, 0, 0, 0, 1, 1, 1, 1, 0, 1,
  0, 1, 1, 0, 0, 0, 0, 1, 1, 0,
  1, 0, 1, 1, 1, 0, 1, 0, 1, 0,
  1, 0, 0, 0, 1, 0, 1, 1, 1, 0,
  1, 0, 1, 0, 1, 0, 1, 1, 1, 0 ;

 Residual =
  0.01463089, 0.008259912, 0.0009736047, 0.005178552, 0.0003064495, 
    0.01201278, 0.003118906, 0.002148788, 0.01049841, 0.0008692471,
  0.003849114, 0.007654977, 0.01492888, 0.002197735, 0.006742722, 
    0.009021605, 0.001459087, 0.004331023, 0.010812, 0.008262091,
  0.01257866, 0.008704971, 0.002768576, 0.009232531, 0.01330433, 0.007751839, 
    0.009392155, 0.007575887, 0.01364494, 0.00619957,
  0.00803203, 0.005139647, 0.001943652, 0.009942327, 0.01403505, 0.009190938, 
    0.01264108, 0.003268627, 0.01354758, 0.0001465497,
  0.003387191, 0.001980827, 0.01361314, 0.01365346, 0.008715869, 0.001312396, 
    0.001753192, 0.01156607, 0.01099193, 0.001306925,
  0.005361948, 0.01159817, 0.001972074, 0.008067487, 0.01132085, 0.004087893, 
    0.008497755, 0.007150275, 0.008349311, 0.006611056,
  0.01040606, 0.01077356, 0.01134574, 0.0005598301, 0.01018253, 0.007158312, 
    0.001502571, 0.009212944, 0.01256872, 0.01100841,
  0.004823484, 0.00101783, 0.0005599536, 0.008386879, 0.00241279, 
    0.004018323, 0.003535679, 0.0002902119, 0.002275296, 0.0005085377,
  0.01472752, 0.00540728, 0.01238197, 0.006183561, 0.003797687, 0.003550663, 
    0.01159673, 0.01006885, 0.01059496, 0.01279733,
  0.007830744, 0.006641545, 0.008306227, 0.009779923, 0.01182831, 0.01338404, 
    0.004636577, 0.002034147, 0.0112639, 0.007902498 ;
}
