netcdf output_1 {
dimensions:
	Scanline = 6 ;
	Field_of_view = 5 ;
	Channel = 22 ;
	Qc_dim = 4 ;
variables:
	short Atm_type(Scanline, Field_of_view) ;
		Atm_type:description = "type of atmosphere:currently missing" ;
		Atm_type:coordinates = "Longitude Latitude" ;
	short BT(Scanline, Field_of_view, Channel) ;
		BT:long_name = "Channel Temperature (K)" ;
		BT:units = "Kelvin" ;
		BT:coordinates = "Longitude Latitude Freq" ;
		BT:scale_factor = 0.01 ;
		BT:_FillValue = -999s ;
		BT:valid_range = 0, 50000 ;
	short CLW(Scanline, Field_of_view) ;
		CLW:long_name = "Cloud liquid Water (mm)" ;
		CLW:units = "mm" ;
		CLW:coordinates = "Longitude Latitude" ;
		CLW:scale_factor = 0.01 ;
		CLW:_FillValue = -999s ;
		CLW:valid_range = 0, 10000 ;
	short ChanSel(Scanline, Field_of_view, Channel) ;
		ChanSel:long_name = "Channels Selection Used in Retrieval" ;
		ChanSel:units = "1" ;
		ChanSel:coordinates = "Longitude Latitude Freq" ;
		ChanSel:_FillValue = -999s ;
		ChanSel:valid_range = 0, 1 ;
	float ChiSqr(Scanline, Field_of_view) ;
		ChiSqr:description = "Convergence rate: <3-good,>10-bad" ;
		ChiSqr:units = "1" ;
		ChiSqr:coordinates = "Longitude Latitude" ;
		ChiSqr:_FillValue = -999.f ;
		ChiSqr:valid_range = 0.f, 1000.f ;
	short CldBase(Scanline, Field_of_view) ;
		CldBase:long_name = "Cloud Base Pressure" ;
		CldBase:scale_factor = 0.1 ;
		CldBase:coordinates = "Longitude Latitude" ;
	short CldThick(Scanline, Field_of_view) ;
		CldThick:long_name = "Cloud Thickness" ;
		CldThick:scale_factor = 0.1 ;
		CldThick:coordinates = "Longitude Latitude" ;
	short CldTop(Scanline, Field_of_view) ;
		CldTop:long_name = "Cloud Top Pressure" ;
		CldTop:scale_factor = 0.1 ;
		CldTop:coordinates = "Longitude Latitude" ;
	short Emis(Scanline, Field_of_view, Channel) ;
		Emis:long_name = "Channel Emissivity" ;
		Emis:units = "1" ;
		Emis:coordinates = "Longitude Latitude Freq" ;
		Emis:scale_factor = 0.0001 ;
		Emis:_FillValue = -999s ;
		Emis:valid_range = 0, 10000 ;
	float Freq(Channel) ;
		Freq:description = "Central Frequencies (GHz)" ;
	short GWP(Scanline, Field_of_view) ;
		GWP:long_name = "Graupel Water Path (mm)" ;
		GWP:units = "mm" ;
		GWP:coordinates = "Longitude Latitude" ;
		GWP:scale_factor = 0.01 ;
		GWP:_FillValue = -999s ;
		GWP:valid_range = 0, 10000 ;
	short IWP(Scanline, Field_of_view) ;
		IWP:long_name = "Ice Water Path (mm)" ;
		IWP:units = "mm" ;
		IWP:coordinates = "Longitude Latitude" ;
		IWP:scale_factor = 0.01 ;
		IWP:_FillValue = -999s ;
		IWP:valid_range = 0, 10000 ;
	short LWP(Scanline, Field_of_view) ;
		LWP:long_name = "Liquid Water Path (mm)" ;
		LWP:units = "mm" ;
		LWP:coordinates = "Longitude Latitude" ;
		LWP:scale_factor = 0.01 ;
		LWP:_FillValue = -999s ;
		LWP:valid_range = 0, 10000 ;
	float LZ_angle(Scanline, Field_of_view) ;
		LZ_angle:long_name = "Local Zenith Angle degree" ;
		LZ_angle:units = "degrees" ;
		LZ_angle:coordinates = "Longitude Latitude" ;
		LZ_angle:_FillValue = -999.f ;
		LZ_angle:valid_range = -70.f, 70.f ;
	float Latitude(Scanline, Field_of_view) ;
		Latitude:long_name = "Latitude of the view (-90,90)" ;
		Latitude:units = "degrees" ;
		Latitude:_FillValue = -999.f ;
		Latitude:valid_range = -90.f, 90.f ;
	float Longitude(Scanline, Field_of_view) ;
		Longitude:long_name = "Longitude of the view (-180,180)" ;
		Longitude:units = "degrees" ;
		Longitude:_FillValue = -999.f ;
		Longitude:valid_range = -180.f, 180.f ;
	short Orb_mode(Scanline) ;
		Orb_mode:description = "0-ascending,1-descending" ;
		Orb_mode:units = "1" ;
		Orb_mode:_FillValue = -999s ;
		Orb_mode:valid_range = 0, 1 ;
	short Polo(Channel) ;
		Polo:description = "Polarizations" ;
	short PrecipType(Scanline, Field_of_view) ;
		PrecipType:long_name = "Precipitation Type (Frozen/Liquid)" ;
		PrecipType:coordinates = "Longitude Latitude" ;
	short Prob_SF(Scanline, Field_of_view) ;
		Prob_SF:long_name = "Probability of falling snow (%)" ;
		Prob_SF:units = "percent" ;
		Prob_SF:coordinates = "Longitude Latitude" ;
		Prob_SF:_FillValue = -999s ;
		Prob_SF:valid_range = 0, 100 ;
	short Qc(Scanline, Field_of_view, Qc_dim) ;
		Qc:description = "Qc: 0-good, 1-usable with problem, 2-bad" ;
	float RAzi_angle(Scanline, Field_of_view) ;
		RAzi_angle:long_name = "Relative Azimuth Angle 0-360 degree" ;
		RAzi_angle:coordinates = "Longitude Latitude" ;
	short RFlag(Scanline, Field_of_view) ;
		RFlag:long_name = "Rain Flag" ;
		RFlag:coordinates = "Longitude Latitude" ;
	short RR(Scanline, Field_of_view) ;
		RR:long_name = "Rain Rate (mm/hr)" ;
		RR:units = "mm/hr" ;
		RR:coordinates = "Longitude Latitude" ;
		RR:scale_factor = 0.1 ;
		RR:_FillValue = -999s ;
		RR:valid_range = 0, 1000 ;
	short RWP(Scanline, Field_of_view) ;
		RWP:long_name = "Rain Water Path (mm)" ;
		RWP:units = "mm" ;
		RWP:coordinates = "Longitude Latitude" ;
		RWP:scale_factor = 0.01 ;
		RWP:_FillValue = -999s ;
		RWP:valid_range = 0, 10000 ;
	short SFR(Scanline, Field_of_view) ;
		SFR:long_name = "Snow Fall Rate in mm/hr" ;
		SFR:units = "mm/hr" ;
		SFR:coordinates = "Longitude Latitude" ;
		SFR:scale_factor = 0.01 ;
		SFR:_FillValue = -999s ;
		SFR:valid_range = 0, 10000 ;
	short SIce(Scanline, Field_of_view) ;
		SIce:long_name = "Sea Ice Concentration (%)" ;
		SIce:units = "percent" ;
		SIce:coordinates = "Longitude Latitude" ;
		SIce:_FillValue = -999s ;
		SIce:valid_range = 0, 100 ;
	short SIce_FY(Scanline, Field_of_view) ;
		SIce_FY:long_name = "First-Year Sea Ice Concentration (%)" ;
		SIce_FY:units = "percent" ;
		SIce_FY:coordinates = "Longitude Latitude" ;
		SIce_FY:_FillValue = -999s ;
		SIce_FY:valid_range = 0, 100 ;
	short SIce_MY(Scanline, Field_of_view) ;
		SIce_MY:long_name = "Multi-Year Sea Ice Concentration (%)" ;
		SIce_MY:units = "percent" ;
		SIce_MY:coordinates = "Longitude Latitude" ;
		SIce_MY:_FillValue = -999s ;
		SIce_MY:valid_range = 0, 100 ;
	short SWE(Scanline, Field_of_view) ;
		SWE:long_name = "Snow Water Equivalent (cm)" ;
		SWE:units = "cm" ;
		SWE:coordinates = "Longitude Latitude" ;
		SWE:scale_factor = 0.01 ;
		SWE:_FillValue = -999s ;
		SWE:valid_range = 0, 10000 ;
	short SWP(Scanline, Field_of_view) ;
		SWP:long_name = "Snow Water Path" ;
		SWP:units = "mm" ;
		SWP:coordinates = "Longitude Latitude" ;
		SWP:scale_factor = 0.01 ;
		SWP:_FillValue = -999s ;
		SWP:valid_range = 0, 10000 ;
	float SZ_angle(Scanline, Field_of_view) ;
		SZ_angle:long_name = "Solar Zenith Angle (-90,90) degree" ;
		SZ_angle:coordinates = "Longitude Latitude" ;
	double ScanTime_UTC(Scanline) ;
		ScanTime_UTC:long_name = "Number of seconds since 00:00:00 UTC" ;
		ScanTime_UTC:units = "seconds" ;
		ScanTime_UTC:_FillValue = -999. ;
		ScanTime_UTC:valid_range = 0., 86400. ;
	short ScanTime_dom(Scanline) ;
		ScanTime_dom:long_name = "Calendar day of the month 1-31" ;
		ScanTime_dom:units = "days" ;
		ScanTime_dom:_FillValue = -999s ;
		ScanTime_dom:valid_range = 1, 31 ;
	short ScanTime_doy(Scanline) ;
		ScanTime_doy:long_name = "julian day 1-366" ;
		ScanTime_doy:units = "days" ;
		ScanTime_doy:_FillValue = -999s ;
		ScanTime_doy:valid_range = 1, 366 ;
	short ScanTime_hour(Scanline) ;
		ScanTime_hour:long_name = "hour of the day 0-23" ;
		ScanTime_hour:units = "hours" ;
		ScanTime_hour:_FillValue = -999s ;
		ScanTime_hour:valid_range = 0, 23 ;
	short ScanTime_minute(Scanline) ;
		ScanTime_minute:long_name = "minute of the hour 0-59" ;
		ScanTime_minute:units = "minutes" ;
		ScanTime_minute:_FillValue = -999s ;
		ScanTime_minute:valid_range = 0, 59 ;
	short ScanTime_month(Scanline) ;
		ScanTime_month:long_name = "Calendar month 1-12" ;
		ScanTime_month:units = "months" ;
		ScanTime_month:_FillValue = -999s ;
		ScanTime_month:valid_range = 1, 12 ;
	short ScanTime_second(Scanline) ;
		ScanTime_second:long_name = "second of the minute 0-59" ;
		ScanTime_second:units = "seconds" ;
		ScanTime_second:_FillValue = -999s ;
		ScanTime_second:valid_range = 0, 59 ;
	short ScanTime_year(Scanline) ;
		ScanTime_year:long_name = "Calendar Year 20XX" ;
		ScanTime_year:units = "years" ;
		ScanTime_year:_FillValue = -999s ;
		ScanTime_year:valid_range = 2011, 2050 ;
	short Sfc_type(Scanline, Field_of_view) ;
		Sfc_type:description = "type of surface:0-ocean,1-sea ice,2-land,3-snow" ;
		Sfc_type:units = "1" ;
		Sfc_type:coordinates = "Longitude Latitude" ;
		Sfc_type:_FillValue = -999s ;
		Sfc_type:valid_range = 0, 3 ;
	short Snow(Scanline, Field_of_view) ;
		Snow:long_name = "Snow Cover" ;
		Snow:units = "1" ;
		Snow:coordinates = "Longitude Latitude" ;
		Snow:_FillValue = -999s ;
		Snow:valid_range = 0, 1 ;
	short SnowGS(Scanline, Field_of_view) ;
		SnowGS:long_name = "Snow Grain Size (mm)" ;
		SnowGS:units = "mm" ;
		SnowGS:coordinates = "Longitude Latitude" ;
		SnowGS:scale_factor = 0.01 ;
		SnowGS:_FillValue = -999s ;
		SnowGS:valid_range = 0, 2000 ;
	short SurfM(Scanline, Field_of_view) ;
		SurfM:long_name = "Surface Moisture" ;
		SurfM:scale_factor = 0.1 ;
		SurfM:coordinates = "Longitude Latitude" ;
	short SurfP(Scanline, Field_of_view) ;
		SurfP:long_name = "Surface Pressure (mb)" ;
		SurfP:units = "millibars" ;
		SurfP:coordinates = "Longitude Latitude" ;
		SurfP:scale_factor = 0.1 ;
		SurfP:_FillValue = -999s ;
		SurfP:valid_range = 0, 12000 ;
	short TPW(Scanline, Field_of_view) ;
		TPW:long_name = "Total Precipitable Water (mm)" ;
		TPW:units = "mm" ;
		TPW:coordinates = "Longitude Latitude" ;
		TPW:scale_factor = 0.1 ;
		TPW:_FillValue = -999s ;
		TPW:valid_range = 0, 2000 ;
	short TSkin(Scanline, Field_of_view) ;
		TSkin:long_name = "Skin Temperature (K)" ;
		TSkin:units = "Kelvin" ;
		TSkin:coordinates = "Longitude Latitude" ;
		TSkin:scale_factor = 0.01 ;
		TSkin:_FillValue = -999s ;
		TSkin:valid_range = 0, 40000 ;
	short WindDir(Scanline, Field_of_view) ;
		WindDir:long_name = "Wind Direction" ;
		WindDir:scale_factor = 0.01 ;
		WindDir:coordinates = "Longitude Latitude" ;
	short WindSp(Scanline, Field_of_view) ;
		WindSp:long_name = "Wind Speed (m/s)" ;
		WindSp:scale_factor = 0.01 ;
		WindSp:coordinates = "Longitude Latitude" ;
	short WindU(Scanline, Field_of_view) ;
		WindU:long_name = "U-direction Wind Speed (m/s)" ;
		WindU:scale_factor = 0.01 ;
		WindU:coordinates = "Longitude Latitude" ;
	short WindV(Scanline, Field_of_view) ;
		WindV:long_name = "V-direction Wind Speed (m/s)" ;
		WindV:scale_factor = 0.01 ;
		WindV:coordinates = "Longitude Latitude" ;
	short YM(Scanline, Field_of_view, Channel) ;
		YM:long_name = "Un-Corrected Channel Temperature (K)" ;
		YM:units = "Kelvin" ;
		YM:coordinates = "Longitude Latitude Freq" ;
		YM:scale_factor = 0.01 ;
		YM:_FillValue = -999s ;
		YM:valid_range = 0, 50000 ;

// global attributes:
		:missing_value = -999 ;
		:notretrievedproduct_value = -888 ;
		:noretrieval_value = -99 ;
		:cdf_version = 4. ;
		:alg_version = 4201 ;
		:dap_version = "v11r4" ;
		:Conventions = "CF-1.5" ;
		:Metadata_Conventions = "CF-1.5, Unidata Dataset Discovery v1.0" ;
		:standard_name_vocabulary = "CF Standard Name Table (version 17, 24 March 2011)" ;
		:project = "Microwave Integrated Retrieval System" ;
		:title = "MIRS IMG" ;
		:summary = "MIRS imaging products including surface emissivity, TPW, CLW, RWP, IWP, LST." ;
		:date_created = "2021-06-30T02:01:08Z" ;
		:institution = "DOC/NOAA/NESDIS/NDE > NPOESS Data Exploitation, NESDIS, NOAA, U.S. Department of Commerce" ;
		:naming_authority = "gov.noaa.nesdis.nde" ;
		:production_site = "NSOF" ;
		:production_environment = "OE" ;
		:satellite_name = "NPP" ;
		:instrument_name = "ATMS" ;
		:creator_name = "DOC/NOAA/NESDIS/STAR > MIRS TEAM, Center for Satellite Applications and Research, NESDIS, NOAA, U.S. Department of Commerce" ;
		:creator_email = "Christopher.Grassotti@noaa.gov, Quanhua.Liu@noaa.gov, Shu-yan.Liu@noaa.gov, ryan.honeyager@noaa.gov, Yong-Keun.Lee@noaa.gov " ;
		:creator_url = "http://www.star.nesdis.noaa.gov/mirs" ;
		:publisher_name = "DOC/NOAA/NESDIS/NDE > NPOESS Data Exploitation, NESDIS, NOAA, U.S. Department of Commerce" ;
		:publisher_email = "NDE_POC@noaa.gov" ;
		:publisher_url = "http://projects.osd.noaa.gov/NDE" ;
		:Metadata_Link = "NDE product-specific output file name" ;
		:references = "http://www.star.nesdis.noaa.gov/mirs/documentation.php" ;
		:history = "Tue Jul 30 17:48:05 2024: ncks -d Scanline,1,12,2 -d Field_of_view,86,94,2 NPR-MIRS-IMG_v11r4_npp_s202106300127066_e202106300127383_c202106300201000.nc output_1.nc\nCreated by MIRS Version 11.4" ;
		:processing_level = "NOAA Level 2 data" ;
		:source = "SATMS_npp_d20210630_t0127066_e0127383_b50120_c20210630015713485030_oebc_ops.h5" ;
		:time_coverage_start = "2021-06-30T01:27:06Z" ;
		:time_coverage_end = "2021-06-30T01:27:38Z" ;
		:cdm_data_type = "Swath" ;
		:geospatial_lat_units = "degrees_north" ;
		:geospatial_lon_units = "degrees_east" ;
		:geospatial_lat_resolution = "100" ;
		:geospatial_lon_resolution = "100" ;
		:geospatial_first_scanline_first_fov_lat = 61.18f ;
		:geospatial_first_scanline_first_fov_lon = 135.75f ;
		:geospatial_first_scanline_last_fov_lat = 69.42f ;
		:geospatial_first_scanline_last_fov_lon = -171.14f ;
		:geospatial_last_scanline_first_fov_lat = 62.38f ;
		:geospatial_last_scanline_first_fov_lon = 133.09f ;
		:geospatial_last_scanline_last_fov_lat = 71.1f ;
		:geospatial_last_scanline_last_fov_lon = -170.7f ;
		:total_number_retrievals = 1152 ;
		:percentage_optimal_retrievals = 0.3125f ;
		:percentage_suboptimal_retrievals = 0.6875f ;
		:percentage_bad_retrievals = 0.f ;
		:start_orbit_number = 50120 ;
		:end_orbit_number = 50120 ;
		:id = "ndepgsl-op-13_2021-06-30T02:01:08Z_0000001764860342_SATMS_npp_d20210630_t0127066_e0127383_b50120_c20210630015713485030_oebc_ops.h5" ;
		:NCO = "netCDF Operators version 5.0.6 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco)" ;
data:

 Atm_type =
  -999, -999, -999, -999, -999,
  -999, -999, -999, -999, -999,
  -999, -999, -999, -999, -999,
  -999, -999, -999, -999, -999,
  -999, -999, -999, -999, -999,
  -999, -999, -999, -999, -999 ;

 BT =
  22327, 22553, 24584, 25405, 25405, 24477, 23433, 23044, 22874, 22877, 
    23030, 23657, 24728, 25747, 26557, 24500, 26503, 26678, 26213, 25708, 
    25076, 24388,
  21454, 21778, 24626, 25336, 25317, 24339, 23404, 22988, 22882, 22870, 
    23110, 23650, 24616, 25911, 26815, 23579, 26248, 26653, 26262, 25888, 
    25060, 24489,
  20583, 20703, 24778, 25420, 25275, 24254, 23307, 22967, 22884, 22926, 
    23216, 23669, 24735, 26131, 27203, 23515, 26303, 26641, 26241, 25768, 
    25210, 24617,
  18802, 18765, 24518, 25360, 25151, 24143, 23200, 22978, 22862, 22898, 
    23093, 23794, 24742, 26033, 26623, 23113, 26509, 26614, 26200, 25725, 
    25061, 24510,
  18595, 18017, 24687, 25325, 25048, 24009, 23120, 22939, 22865, 22946, 
    23224, 23879, 24829, 26147, 27059, 22539, 26383, 26362, 25866, 25253, 
    24545, 23854,
  20793, 21116, 23628, 24840, 25233, 24424, 23390, 23045, 22901, 22904, 
    23094, 23688, 24648, 25831, 26676, 22575, 25726, 26585, 26195, 25717, 
    25064, 24363,
  21377, 21586, 24734, 25380, 25331, 24369, 23401, 23045, 22868, 22934, 
    23189, 23708, 24567, 25960, 26841, 23692, 26248, 26683, 26257, 25791, 
    25193, 24557,
  21381, 21420, 25117, 25561, 25226, 24274, 23292, 22993, 22911, 22893, 
    23138, 23665, 24838, 26055, 26847, 24056, 26334, 26585, 26140, 25814, 
    25120, 24504,
  19667, 19643, 24743, 25396, 25127, 24148, 23195, 22934, 22871, 22917, 
    23140, 23828, 24779, 26136, 27013, 23313, 26553, 26566, 26085, 25653, 
    25054, 24377,
  18796, 18249, 24810, 25396, 25050, 24028, 23159, 22958, 22904, 22927, 
    23254, 23769, 24910, 26096, 27232, 22485, 26377, 26435, 25985, 25404, 
    24735, 24056,
  20498, 20619, 24167, 25066, 25273, 24456, 23441, 23055, 22845, 22994, 
    23204, 23619, 24720, 25987, 26769, 23008, 26075, 26562, 26192, 25755, 
    25061, 24573,
  21974, 22034, 24987, 25431, 25308, 24348, 23367, 23050, 22914, 22895, 
    23120, 23721, 24623, 25823, 26791, 23833, 26149, 26594, 26254, 25766, 
    25196, 24606,
  22286, 22455, 25270, 25612, 25241, 24266, 23347, 23022, 22882, 23061, 
    23197, 23677, 24769, 25901, 26953, 24352, 26322, 26612, 26150, 25802, 
    25136, 24695,
  20622, 20769, 25003, 25495, 25182, 24147, 23257, 23022, 22900, 23025, 
    23304, 23842, 24848, 26110, 26759, 23649, 26478, 26571, 26192, 25728, 
    25063, 24466,
  19327, 18919, 25100, 25537, 25062, 24009, 23201, 22992, 22929, 23026, 
    23256, 23809, 24836, 26290, 27335, 23116, 26365, 26440, 25947, 25510, 
    24884, 24272,
  21249, 21254, 24759, 25349, 25313, 24440, 23466, 23067, 22965, 23009, 
    23255, 23621, 24619, 25850, 27194, 24105, 26399, 26501, 26057, 25603, 
    24990, 24414,
  22658, 22722, 24961, 25453, 25265, 24357, 23360, 23024, 22940, 23014, 
    23245, 23711, 24671, 25754, 27012, 23734, 26119, 26526, 26154, 25713, 
    25146, 24615,
  22959, 23177, 25363, 25634, 25235, 24239, 23334, 23023, 22907, 23019, 
    23186, 23742, 24777, 26127, 26904, 24337, 26303, 26572, 26112, 25707, 
    25029, 24396,
  21486, 21662, 25154, 25560, 25188, 24203, 23268, 23049, 22949, 23043, 
    23274, 23804, 24848, 26228, 27015, 24075, 26566, 26510, 26126, 25620, 
    24987, 24489,
  19966, 19685, 25024, 25462, 25036, 24029, 23177, 23025, 22970, 23030, 
    23250, 23833, 24928, 26123, 26876, 23233, 26472, 26459, 26075, 25576, 
    25050, 24462,
  22101, 22142, 24626, 25300, 25300, 24421, 23492, 23108, 22989, 22996, 
    23273, 23624, 24619, 26074, 26893, 23896, 26110, 26501, 26128, 25586, 
    25049, 24481,
  22985, 23104, 25074, 25606, 25321, 24344, 23442, 23067, 22944, 22979, 
    23243, 23825, 24698, 26006, 27066, 24230, 26434, 26519, 26068, 25716, 
    25108, 24535,
  23325, 23451, 25676, 25810, 25325, 24232, 23370, 23076, 22937, 23023, 
    23175, 23773, 24758, 26123, 26956, 25236, 26625, 26515, 26135, 25720, 
    25029, 24403,
  22237, 22340, 25362, 25622, 25147, 24160, 23253, 23042, 22990, 22986, 
    23282, 23852, 24876, 26304, 27106, 24686, 26632, 26416, 25971, 25497, 
    24880, 24287,
  20683, 20418, 24990, 25420, 25000, 24034, 23200, 23015, 22971, 23025, 
    23331, 23892, 24923, 26416, 26846, 23170, 26333, 26315, 25872, 25491, 
    24835, 24308,
  22590, 22687, 24808, 25303, 25314, 24410, 23474, 23116, 22966, 23030, 
    23196, 23638, 24636, 25891, 26881, 24034, 26215, 26377, 25982, 25584, 
    24962, 24423,
  23025, 23150, 25193, 25587, 25349, 24383, 23407, 23090, 22970, 22979, 
    23231, 23757, 24766, 26025, 26894, 24597, 26450, 26373, 25997, 25490, 
    24876, 24390,
  23403, 23510, 25850, 25891, 25304, 24246, 23363, 23124, 22967, 23032, 
    23266, 23794, 24782, 26245, 26928, 25768, 26897, 26420, 25934, 25489, 
    24899, 24318,
  22797, 22937, 25424, 25596, 25175, 24149, 23293, 23056, 22994, 23090, 
    23257, 23835, 24904, 25935, 27034, 24841, 26579, 26436, 25983, 25501, 
    24902, 24358,
  21439, 21265, 25131, 25468, 25006, 23978, 23199, 23067, 23015, 23028, 
    23336, 23936, 24811, 26224, 27077, 23546, 26454, 26276, 25912, 25458, 
    24844, 24264 ;

 CLW =
  4, 0, 0, 2, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 2, 7, 5, 0 ;

 ChanSel =
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1 ;

 ChiSqr =
  0.3278425, 0.1270331, 0.5191541, 0.1502331, 0.1583424,
  0.2056985, 0.09662999, 0.4452049, 0.1618346, 0.2081715,
  0.7202161, 0.7179015, 0.3983652, 0.2625816, 0.9757569,
  0.264237, 0.8345357, 0.2943406, 0.1115318, 0.5097764,
  0.169713, 0.409044, 0.1654734, 0.1077542, 0.3691869,
  0.6970016, 0.4721045, 0.4847079, 0.4702559, 0.4022827 ;

 CldBase =
  -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888 ;

 CldThick =
  -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888 ;

 CldTop =
  -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888 ;

 Emis =
  7664, 7844, 7419, 7437, 7450, 7460, 7470, 7477, 7483, 7503, 7503, 7503, 
    7503, 7503, 7503, 8176, 8189, 8189, 8189, 8189, 8189, 8189,
  7207, 7421, 7496, 7509, 7519, 7526, 7533, 7537, 7542, 7557, 7557, 7557, 
    7557, 7557, 7557, 7808, 8056, 8056, 8056, 8056, 8056, 8056,
  6756, 7105, 7499, 7507, 7513, 7517, 7522, 7524, 7527, 7535, 7535, 7535, 
    7535, 7535, 7535, 7803, 7831, 7831, 7831, 7831, 7831, 7831,
  5775, 6024, 6681, 6711, 6732, 6748, 6764, 6774, 6785, 6819, 6819, 6819, 
    6819, 6819, 6819, 7102, 7947, 8063, 8063, 8063, 8063, 8063,
  5670, 5923, 6789, 6820, 6841, 6857, 6873, 6883, 6895, 6928, 6928, 6928, 
    6928, 6928, 6928, 7000, 8029, 8141, 8141, 8141, 8141, 8141,
  7151, 7229, 6826, 6859, 6882, 6899, 6916, 6927, 6939, 6975, 6975, 6975, 
    6975, 6975, 6975, 7525, 8182, 8182, 8182, 8182, 8182, 8182,
  7152, 7402, 7560, 7571, 7579, 7584, 7590, 7593, 7597, 7609, 7609, 7609, 
    7609, 7609, 7609, 7851, 8010, 8010, 8010, 8010, 8010, 8010,
  7142, 7510, 7958, 7957, 7956, 7955, 7955, 7954, 7953, 7952, 7952, 7952, 
    7952, 7952, 7952, 8116, 7899, 7898, 7898, 7898, 7899, 7899,
  6216, 6461, 7131, 7159, 7178, 7193, 7207, 7217, 7227, 7258, 7258, 7258, 
    7258, 7258, 7258, 7452, 8253, 8358, 8358, 8358, 8358, 8358,
  5806, 6037, 6985, 7012, 7032, 7046, 7060, 7069, 7080, 7111, 7111, 7111, 
    7111, 7111, 7111, 7010, 8103, 8208, 8208, 8208, 8208, 8208,
  6895, 7148, 7235, 7256, 7270, 7281, 7291, 7298, 7305, 7328, 7328, 7328, 
    7328, 7328, 7328, 7765, 8086, 8086, 8086, 8086, 8086, 8086,
  7574, 7861, 8078, 8077, 8077, 8077, 8077, 8076, 8076, 8075, 8075, 8075, 
    8075, 8075, 8075, 8248, 8048, 8048, 8048, 8048, 8048, 8049,
  7592, 7901, 8200, 8197, 8194, 8192, 8190, 8188, 8187, 8183, 8183, 8183, 
    8183, 8183, 8183, 8303, 8039, 8039, 8039, 8039, 8039, 8039,
  6567, 6941, 7499, 7501, 7503, 7504, 7504, 7505, 7505, 7507, 7507, 7507, 
    7507, 7507, 7507, 7602, 7570, 7570, 7570, 7570, 7570, 7570,
  5890, 6418, 7360, 7359, 7359, 7358, 7357, 7357, 7356, 7355, 7355, 7355, 
    7355, 7355, 7355, 7486, 7309, 7309, 7309, 7309, 7309, 7310,
  7080, 7410, 7679, 7692, 7701, 7708, 7714, 7718, 7723, 7737, 7737, 7737, 
    7737, 7737, 7737, 8135, 8209, 8209, 8209, 8209, 8209, 8209,
  7903, 8112, 8143, 8142, 8141, 8140, 8140, 8139, 8138, 8137, 8137, 8137, 
    8137, 8137, 8137, 8257, 8082, 8081, 8081, 8082, 8082, 8082,
  7913, 8168, 8362, 8354, 8349, 8345, 8341, 8338, 8335, 8326, 8326, 8326, 
    8326, 8326, 8326, 8344, 8036, 8036, 8036, 8036, 8036, 8036,
  6944, 7284, 7726, 7726, 7726, 7726, 7726, 7725, 7725, 7725, 7725, 7725, 
    7725, 7725, 7725, 7821, 7720, 7720, 7720, 7720, 7720, 7720,
  6145, 6574, 7317, 7317, 7317, 7316, 7316, 7315, 7315, 7315, 7315, 7315, 
    7315, 7315, 7315, 7356, 7295, 7295, 7295, 7295, 7296, 7296,
  7584, 7766, 7681, 7696, 7706, 7713, 7720, 7724, 7729, 7745, 7745, 7745, 
    7745, 7745, 7745, 8074, 8262, 8262, 8262, 8262, 8262, 8262,
  7987, 8130, 8038, 8046, 8052, 8056, 8062, 8065, 8068, 8077, 8077, 8077, 
    8077, 8077, 8077, 8367, 8397, 8397, 8397, 8397, 8397, 8397,
  7878, 8192, 8503, 8494, 8487, 8482, 8477, 8474, 8470, 8460, 8460, 8460, 
    8460, 8460, 8460, 8519, 8101, 8101, 8101, 8101, 8101, 8101,
  7298, 7641, 8057, 8054, 8052, 8050, 8048, 8047, 8045, 8042, 8042, 8042, 
    8042, 8042, 8042, 8144, 7915, 7915, 7915, 7915, 7915, 7915,
  6567, 6916, 7470, 7467, 7465, 7463, 7462, 7460, 7459, 7455, 7455, 7455, 
    7455, 7455, 7455, 7416, 7333, 7333, 7333, 7333, 7333, 7333,
  7840, 8059, 8034, 8041, 8045, 8049, 8052, 8054, 8056, 8064, 8064, 8064, 
    8064, 8064, 8064, 8365, 8304, 8303, 8303, 8304, 8304, 8304,
  7912, 8034, 8095, 8105, 8113, 8118, 8124, 8127, 8132, 8143, 8143, 8143, 
    8143, 8143, 8143, 8442, 8605, 8681, 8681, 8681, 8681, 8681,
  7838, 8000, 8345, 8351, 8356, 8359, 8364, 8366, 8368, 8376, 8376, 8376, 
    8376, 8376, 8376, 8510, 8633, 8633, 8633, 8633, 8633, 8633,
  7797, 7948, 8188, 8201, 8210, 8217, 8224, 8228, 8234, 8249, 8249, 8249, 
    8249, 8249, 8249, 8445, 8750, 8825, 8825, 8825, 8825, 8825,
  6896, 7206, 7683, 7675, 7670, 7666, 7662, 7659, 7657, 7648, 7648, 7648, 
    7648, 7648, 7648, 7528, 7365, 7365, 7365, 7365, 7365, 7365 ;

 Freq = 23.8, 31.4, 50.3, 51.76, 52.8, 53.596, 54.4, 54.94, 55.5, 57.29, 
    57.29, 57.29, 57.29, 57.29, 57.29, 88.2, 165.5, 183.31, 183.31, 183.31, 
    183.31, 183.31 ;

 GWP =
  0, _, _, _, _,
  _, _, _, _, _,
  _, _, _, _, _,
  _, _, _, _, _,
  _, 0, _, _, _,
  _, _, 0, _, _ ;

 IWP =
  _, _, _, _, _,
  _, _, _, _, _,
  _, _, _, _, _,
  _, _, _, _, _,
  _, _, _, _, _,
  _, _, _, _, _ ;

 LWP =
  4, -998, -998, -998, -998,
  -998, -998, -998, -998, -998,
  -998, -998, -998, -998, -998,
  -998, -998, -998, -998, -998,
  -998, 0, -998, -998, -998,
  -998, -998, 7, -998, -998 ;

 LZ_angle =
  50.15001, 53.07, 56.06001, 59.21, 62.46,
  50.15001, 53.07, 56.08001, 59.18999, 62.47999,
  50.16999, 53.05, 56.09, 59.18999, 62.46998,
  50.16999, 53.08001, 56.08001, 59.21, 62.45,
  50.15001, 53.08001, 56.07, 59.2, 62.47999,
  50.15999, 53.07, 56.09, 59.18001, 62.48999 ;

 Latitude =
  69.59, 69.64, 69.67, 69.67, 69.62,
  69.9, 69.95, 69.98, 69.98, 69.93,
  70.21, 70.26, 70.29, 70.29, 70.24,
  70.52, 70.57, 70.6, 70.6, 70.55,
  70.83, 70.88, 70.91, 70.91, 70.85,
  71.14, 71.2, 71.23, 71.22, 71.16 ;

 Longitude =
  177.29, 179.29, -178.47, -175.86, -172.85,
  177.19, 179.21, -178.5, -175.88, -172.78,
  177.1, 179.13, -178.52, -175.87, -172.75,
  177, 179.07, -178.57, -175.85, -172.71,
  176.88, 179, -178.61, -175.85, -172.63,
  176.78, 178.92, -178.63, -175.86, -172.56 ;

 Orb_mode = 0, 0, 0, 0, 0, 0 ;

 Polo = 2, 2, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 2, 3, 3, 3, 3, 3, 3 ;

 PrecipType =
  -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888 ;

 Prob_SF =
  _, _, _, _, _,
  _, _, _, _, _,
  _, _, _, _, _,
  _, _, _, _, _,
  _, _, _, _, _,
  _, _, _, _, _ ;

 Qc =
  0, 0, 160, 8192,
  0, 0, 128, 0,
  0, 0, 128, 0,
  0, 0, 32, 4096,
  0, 0, 0, 4096,
  0, 0, 128, 0,
  0, 0, 128, 0,
  0, 0, 128, 0,
  0, 0, 0, 4096,
  0, 0, 0, 4096,
  0, 0, 128, 0,
  0, 0, 128, 0,
  0, 0, 128, 0,
  0, 0, 128, 0,
  0, 0, 128, 0,
  0, 0, 128, 0,
  0, 0, 128, 0,
  0, 0, 128, 0,
  0, 0, 128, 0,
  0, 0, 128, 0,
  0, 0, 128, 0,
  0, 0, 128, 8192,
  0, 0, 128, 0,
  0, 0, 128, 0,
  0, 0, 128, 0,
  1, 0, 144, 0,
  0, 0, 32, 4096,
  0, 0, 160, 8192,
  0, 0, 32, 4096,
  1, 0, 144, 0 ;

 RAzi_angle =
  -95.03, -93.16, -91.06, -88.61, -85.79,
  -95.07, -93.17, -91.02, -88.56, -85.65,
  -95.09, -93.18, -90.97, -88.48, -85.54,
  -95.12, -93.17, -90.95, -88.38, -85.42,
  -95.18, -93.17, -90.92, -88.3, -85.27,
  -95.21, -93.18, -90.86, -88.25, -85.12 ;

 RFlag =
  -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888 ;

 RR =
  0, _, _, _, _,
  _, _, _, _, _,
  _, _, _, _, _,
  _, _, _, _, _,
  _, 0, _, _, _,
  _, _, 0, _, _ ;

 RWP =
  0, _, _, _, _,
  _, _, _, _, _,
  _, _, _, _, _,
  _, _, _, _, _,
  _, 0, _, _, _,
  _, _, 0, _, _ ;

 SFR =
  _, _, _, _, _,
  _, _, _, _, _,
  _, _, _, _, _,
  _, _, _, _, _,
  _, _, _, _, _,
  _, _, _, _, _ ;

 SIce =
  _, 58, 52, 0, 0,
  52, 58, 62, 38, 0,
  52, 70, 72, 0, 0,
  60, 76, 78, 56, 0,
  68, _, 80, 66, 46,
  76, 76, _, 76, 0 ;

 SIce_FY =
  _, 58, 52, 0, 0,
  52, 58, 62, 38, 0,
  52, 70, 72, 0, 0,
  60, 76, 78, 56, 0,
  68, _, 80, 66, 45,
  76, 76, _, 76, 0 ;

 SIce_MY =
  _, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, _, 0, 0, 0,
  0, 0, _, 0, 0 ;

 SWE =
  0, _, _, _, _,
  _, _, _, _, _,
  _, _, _, _, _,
  _, _, _, _, _,
  _, 0, _, _, _,
  _, _, 0, _, _ ;

 SWP =
  _, _, _, _, _,
  _, _, _, _, _,
  _, _, _, _, _,
  _, _, _, _, _,
  _, _, _, _, _,
  _, _, _, _, _ ;

 SZ_angle =
  47.68, 48.01, 48.39, 48.83, 49.36,
  47.95, 48.28, 48.66, 49.1, 49.63,
  48.23, 48.56, 48.93, 49.37, 49.9,
  48.51, 48.83, 49.21, 49.64, 50.16,
  48.78, 49.11, 49.48, 49.91, 50.43,
  49.06, 49.38, 49.76, 50.18, 50.7 ;

 ScanTime_UTC = 5229.00048828125, 5234.00048828125, 5240.00048828125, 
    5245.00048828125, 5250.00048828125, 5256.00048828125 ;

 ScanTime_dom = 30, 30, 30, 30, 30, 30 ;

 ScanTime_doy = 181, 181, 181, 181, 181, 181 ;

 ScanTime_hour = 1, 1, 1, 1, 1, 1 ;

 ScanTime_minute = 27, 27, 27, 27, 27, 27 ;

 ScanTime_month = 6, 6, 6, 6, 6, 6 ;

 ScanTime_second = 9, 14, 20, 25, 30, 36 ;

 ScanTime_year = 2021, 2021, 2021, 2021, 2021, 2021 ;

 Sfc_type =
  2, 1, 1, 0, 0,
  1, 1, 1, 1, 0,
  1, 1, 1, 0, 0,
  1, 1, 1, 1, 0,
  1, 2, 1, 1, 1,
  1, 1, 2, 1, 0 ;

 Snow =
  0, _, _, _, _,
  _, _, _, _, _,
  _, _, _, _, _,
  _, _, _, _, _,
  _, 0, _, _, _,
  _, _, 0, _, _ ;

 SnowGS =
  0, _, _, _, _,
  _, _, _, _, _,
  _, _, _, _, _,
  _, _, _, _, _,
  _, 0, _, _, _,
  _, _, 0, _, _ ;

 SurfM =
  -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888 ;

 SurfP =
  10046, 9930, 9930, 9930, 9930,
  9930, 9930, 9930, 9930, 9930,
  9930, 9930, 9930, 9930, 9930,
  9930, 9930, 9930, 9930, 9930,
  9930, 10092, 9930, 9930, 9930,
  9930, 10084, 9796, 10084, 9930 ;

 TPW =
  109, 107, 108, 103, 101,
  89, 107, 110, 106, 96,
  111, 106, 108, 123, 116,
  122, 110, 108, 130, 123,
  103, 119, 128, 133, 124,
  126, 110, 124, 95, 130 ;

 TSkin =
  27460, 27593, 27982, 27901, 27718,
  27122, 27666, 27847, 27840, 27733,
  27385, 27513, 27718, 28090, 28389,
  27715, 27420, 27685, 27993, 28310,
  27460, 27463, 27945, 27978, 27967,
  27305, 27795, 28165, 27668, 28025 ;

 WindDir =
  -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888 ;

 WindSp =
  -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888 ;

 WindU =
  -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888 ;

 WindV =
  -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888 ;

 YM =
  22619, 22707, 24720, 25360, 25272, 24389, 23362, 22925, 22768, 22824, 
    22970, 23608, 24653, 25651, 26487, 24562, 26332, 26521, 26087, 25591, 
    24965, 24324,
  21757, 21949, 24710, 25252, 25172, 24250, 23328, 22866, 22775, 22816, 
    23047, 23598, 24539, 25816, 26741, 23607, 26072, 26493, 26135, 25772, 
    24947, 24425,
  20878, 20881, 24797, 25290, 25118, 24163, 23227, 22841, 22775, 22870, 
    23150, 23614, 24653, 26029, 27129, 23483, 26110, 26471, 26109, 25648, 
    25094, 24552,
  19142, 19003, 24470, 25177, 24984, 24043, 23117, 22850, 22750, 22842, 
    23026, 23736, 24656, 25926, 26548, 23016, 26297, 26435, 26060, 25604, 
    24942, 24440,
  19011, 18355, 24562, 25105, 24873, 23904, 23031, 22809, 22753, 22889, 
    23157, 23818, 24738, 26038, 26982, 22368, 26160, 26176, 25724, 25128, 
    24421, 23778,
  21085, 21270, 23764, 24795, 25100, 24336, 23319, 22926, 22795, 22851, 
    23034, 23639, 24573, 25735, 26606, 22637, 25556, 26428, 26069, 25600, 
    24952, 24299,
  21680, 21757, 24818, 25296, 25186, 24280, 23326, 22923, 22761, 22880, 
    23126, 23656, 24490, 25865, 26768, 23720, 26072, 26523, 26131, 25675, 
    25080, 24493,
  21676, 21598, 25136, 25431, 25069, 24183, 23212, 22868, 22802, 22837, 
    23072, 23610, 24756, 25954, 26773, 24024, 26141, 26415, 26007, 25694, 
    25004, 24440,
  20007, 19881, 24695, 25213, 24960, 24048, 23112, 22806, 22759, 22861, 
    23073, 23770, 24693, 26029, 26938, 23216, 26341, 26387, 25946, 25533, 
    24935, 24307,
  19212, 18587, 24685, 25176, 24875, 23923, 23070, 22828, 22792, 22870, 
    23187, 23707, 24819, 25987, 27156, 22314, 26154, 26250, 25843, 25279, 
    24611, 23980,
  20790, 20773, 24303, 25021, 25140, 24368, 23370, 22936, 22739, 22941, 
    23144, 23570, 24645, 25891, 26698, 23070, 25904, 26404, 26066, 25638, 
    24949, 24509,
  22277, 22205, 25071, 25347, 25163, 24259, 23291, 22928, 22807, 22841, 
    23057, 23669, 24546, 25728, 26717, 23861, 25973, 26434, 26128, 25650, 
    25083, 24542,
  22581, 22633, 25289, 25482, 25084, 24175, 23267, 22896, 22773, 23005, 
    23131, 23622, 24687, 25800, 26879, 24320, 26129, 26442, 26018, 25682, 
    25020, 24630,
  20962, 21007, 24955, 25312, 25015, 24047, 23174, 22894, 22788, 22969, 
    23237, 23784, 24762, 26003, 26684, 23552, 26266, 26392, 26053, 25607, 
    24944, 24396,
  19743, 19257, 24975, 25318, 24887, 23904, 23112, 22862, 22818, 22969, 
    23189, 23747, 24745, 26181, 27259, 22945, 26142, 26254, 25804, 25385, 
    24760, 24196,
  21541, 21408, 24895, 25304, 25180, 24352, 23395, 22948, 22859, 22956, 
    23195, 23572, 24544, 25754, 27123, 24167, 26228, 26344, 25931, 25486, 
    24879, 24350,
  22961, 22893, 25045, 25369, 25120, 24268, 23284, 22902, 22833, 22960, 
    23182, 23659, 24594, 25659, 26938, 23762, 25943, 26366, 26028, 25598, 
    25033, 24551,
  23254, 23355, 25382, 25504, 25078, 24148, 23254, 22897, 22798, 22963, 
    23120, 23687, 24695, 26026, 26831, 24305, 26110, 26401, 25979, 25587, 
    24913, 24331,
  21826, 21900, 25106, 25377, 25021, 24103, 23185, 22921, 22837, 22987, 
    23206, 23746, 24762, 26121, 26940, 23978, 26354, 26331, 25987, 25500, 
    24868, 24419,
  20382, 20023, 24899, 25243, 24861, 23924, 23088, 22895, 22858, 22973, 
    23183, 23771, 24837, 26014, 26800, 23062, 26249, 26273, 25932, 25451, 
    24926, 24386,
  22393, 22296, 24762, 25255, 25167, 24333, 23421, 22989, 22883, 22943, 
    23213, 23575, 24544, 25978, 26822, 23958, 25940, 26344, 26001, 25469, 
    24937, 24417,
  23288, 23275, 25158, 25522, 25176, 24255, 23366, 22945, 22837, 22926, 
    23180, 23773, 24621, 25910, 26992, 24258, 26257, 26359, 25941, 25600, 
    24995, 24471,
  23620, 23629, 25695, 25681, 25168, 24141, 23290, 22951, 22829, 22967, 
    23109, 23718, 24676, 26022, 26882, 25204, 26432, 26345, 26003, 25600, 
    24913, 24338,
  22577, 22578, 25315, 25439, 24980, 24060, 23170, 22914, 22879, 22930, 
    23215, 23794, 24790, 26197, 27031, 24589, 26420, 26237, 25832, 25377, 
    24761, 24218,
  21099, 20756, 24865, 25200, 24825, 23929, 23111, 22885, 22859, 22968, 
    23264, 23830, 24832, 26307, 26770, 22999, 26110, 26129, 25729, 25366, 
    24711, 24232,
  22882, 22841, 24944, 25258, 25181, 24322, 23403, 22997, 22860, 22977, 
    23136, 23589, 24561, 25795, 26810, 24096, 26044, 26220, 25856, 25467, 
    24851, 24359,
  23328, 23321, 25277, 25503, 25204, 24294, 23331, 22968, 22863, 22926, 
    23168, 23705, 24689, 25929, 26821, 24625, 26274, 26213, 25870, 25374, 
    24763, 24326,
  23698, 23688, 25869, 25762, 25147, 24155, 23283, 22998, 22858, 22976, 
    23200, 23739, 24700, 26144, 26854, 25735, 26704, 26250, 25801, 25369, 
    24783, 24253,
  23137, 23175, 25376, 25413, 25008, 24049, 23210, 22928, 22882, 23034, 
    23189, 23777, 24818, 25828, 26959, 24744, 26368, 26257, 25844, 25381, 
    24783, 24288,
  21855, 21603, 25006, 25248, 24831, 23873, 23110, 22937, 22903, 22971, 
    23269, 23874, 24720, 26115, 27001, 23375, 26231, 26091, 25769, 25333, 
    24720, 24188 ;
}
