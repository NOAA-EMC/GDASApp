netcdf sss_smos_1_sub {
dimensions:
	n_grid_points = 52 ;
variables:
	short Dg_quality_SSS_corr(n_grid_points) ;
		Dg_quality_SSS_corr:_FillValue = 999US ;
		string Dg_quality_SSS_corr:_Unsigned = "true" ;
	float Latitude(n_grid_points) ;
		string Latitude:units = "deg" ;
		Latitude:_FillValue = -999.f ;
	float Longitude(n_grid_points) ;
		string Longitude:units = "deg" ;
		Longitude:_FillValue = -999.f ;
	float Mean_acq_time(n_grid_points) ;
		string Mean_acq_time:units = "dd" ;
		Mean_acq_time:_FillValue = -999.f ;
	float SSS_corr(n_grid_points) ;
		string SSS_corr:units = "psu" ;
		SSS_corr:_FillValue = -999.f ;
	float Sigma_SSS_corr(n_grid_points) ;
		string Sigma_SSS_corr:units = "psu" ;
		Sigma_SSS_corr:_FillValue = -999.f ;

// global attributes:
		string :creation_date = "UTC=2021-07-01T03:51:46" ;
		string :total_number_of_grid_points = "106350" ;
		string :FH\:File_Name = "SM_OPER_MIR_OSUDP2_20210630T210913_20210630T220228_700_001_1" ;
		string :FH\:File_Description = "L2 Ocean Salinity Output User Data Product." ;
		string :FH\:Notes = "The UDP (User Data Product) is designed for oceanographics and high level centers, it includes geophysical parameters, a theoretical estimate of their accuracy, flags and descriptors of the product quality." ;
		string :FH\:Mission = "SMOS" ;
		string :FH\:File_Class = "OPER" ;
		string :FH\:File_Type = "MIR_OSUDP2" ;
		string :FH\:File_Version = "0001" ;
		string :FH\:Validity_Period\:Validity_Start = "UTC=2021-06-30T21:09:13" ;
		string :FH\:Validity_Period\:Validity_Stop = "UTC=2021-06-30T22:02:28" ;
		string :FH\:Source\:System = "DPGS" ;
		string :FH\:Source\:Creator = "L2OP" ;
		string :FH\:Source\:Creator_Version = "700" ;
		string :FH\:Source\:Creation_Date = "UTC=2021-07-01T03:44:36" ;
		string :VH\:SPH\:QI\:Total_Selected_L1c_Grid_Points = "80650" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:Retrieval_Scheme = "1" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:Land_Rejected = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:Too_Close_To_Land_Rejected = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:Ice_Rejected = "9107" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:Missing_ECMWF_Rejected = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:Too_Few_Measurements_Rejected = "14105" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:Good_Quality_Grid_Points = "49030" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:Poor_Quality_Grid_Points = "10594" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:SQ\:Grid_Point_Type = "Sea" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:SQ\:SSS_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:SQ\:SST_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:SQ\:WS_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:SQ\:Good_Quality = "42416" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:SQ\:Good_Quality_Retrieved = "33881" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:SQ\:Good_Quality_Retrieved_Average_Sigma = "1.300973" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:SQ\:Good_Quality_Failed_Outside_Valid_Range = "138" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:SQ\:Good_Quality_Failed_Sigma_Too_High = "456" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:SQ\:Good_Quality_Failed_Poor_Fit = "7974" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:SQ\:Good_Quality_Failed_Marquardt = "50" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:SQ\:Good_Quality_Failed_Maxiter = "489" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:SQ\:Good_Quality_Failed_OOLUT = "549" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:SQ\:Poor_Quality = "7258" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:SQ\:Poor_Quality_Retrieved = "5481" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:SQ\:Poor_Quality_Retrieved_Average_Sigma = "2.500925" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:NCQ\:Grid_Point_Type = "Near_Coast" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:NCQ\:SSS_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:NCQ\:SST_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:NCQ\:WS_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:NCQ\:Good_Quality = "6614" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:NCQ\:Good_Quality_Retrieved = "3994" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:NCQ\:Good_Quality_Retrieved_Average_Sigma = "2.145041" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:NCQ\:Good_Quality_Failed_Outside_Valid_Range = "331" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:NCQ\:Good_Quality_Failed_Sigma_Too_High = "780" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:NCQ\:Good_Quality_Failed_Poor_Fit = "2270" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:NCQ\:Good_Quality_Failed_Marquardt = "175" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:NCQ\:Good_Quality_Failed_Maxiter = "307" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:NCQ\:Good_Quality_Failed_OOLUT = "993" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:NCQ\:Poor_Quality = "3336" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:NCQ\:Poor_Quality_Retrieved = "2402" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:NCQ\:Poor_Quality_Retrieved_Average_Sigma = "2.491391" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_0\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_0\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_0\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_0\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_0\:Good_Quality = "40" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_0\:Good_Quality_Retrieved = "13" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_0\:Good_Quality_Retrieved_Average_Sigma = "2.271775" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_0\:Good_Quality_Failed_Outside_Valid_Range = "11" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_0\:Good_Quality_Failed_Sigma_Too_High = "13" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_0\:Good_Quality_Failed_Poor_Fit = "26" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_0\:Good_Quality_Failed_Marquardt = "6" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_0\:Good_Quality_Failed_Maxiter = "6" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_0\:Good_Quality_Failed_OOLUT = "14" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_0\:Poor_Quality = "11" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_0\:Poor_Quality_Retrieved = "6" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_0\:Poor_Quality_Retrieved_Average_Sigma = "4.644665" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_1\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_1\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_1\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_1\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_1\:Good_Quality = "32" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_1\:Good_Quality_Retrieved = "25" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_1\:Good_Quality_Retrieved_Average_Sigma = "2.331885" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_1\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_1\:Good_Quality_Failed_Sigma_Too_High = "3" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_1\:Good_Quality_Failed_Poor_Fit = "6" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_1\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_1\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_1\:Good_Quality_Failed_OOLUT = "4" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_1\:Poor_Quality = "185" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_1\:Poor_Quality_Retrieved = "8" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_1\:Poor_Quality_Retrieved_Average_Sigma = "4.768177" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_2\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_2\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_2\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_2\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_2\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_2\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_2\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_2\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_2\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_2\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_2\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_2\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_2\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_2\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_2\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_2\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_3\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_3\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_3\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_3\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_3\:Good_Quality = "6" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_3\:Good_Quality_Retrieved = "6" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_3\:Good_Quality_Retrieved_Average_Sigma = "1.849856" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_3\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_3\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_3\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_3\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_3\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_3\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_3\:Poor_Quality = "92" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_3\:Poor_Quality_Retrieved = "61" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_3\:Poor_Quality_Retrieved_Average_Sigma = "3.938132" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_4\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_4\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_4\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_4\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_4\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_4\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_4\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_4\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_4\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_4\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_4\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_4\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_4\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_4\:Poor_Quality = "371" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_4\:Poor_Quality_Retrieved = "214" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_4\:Poor_Quality_Retrieved_Average_Sigma = "4.211347" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_5\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_5\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_5\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_5\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_5\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_5\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_5\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_5\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_5\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_5\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_5\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_5\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_5\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_5\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_5\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_5\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_6\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_6\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_6\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_6\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_6\:Good_Quality = "127" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_6\:Good_Quality_Retrieved = "36" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_6\:Good_Quality_Retrieved_Average_Sigma = "0.556612" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_6\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_6\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_6\:Good_Quality_Failed_Poor_Fit = "87" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_6\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_6\:Good_Quality_Failed_Maxiter = "9" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_6\:Good_Quality_Failed_OOLUT = "16" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_6\:Poor_Quality = "16" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_6\:Poor_Quality_Retrieved = "9" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_6\:Poor_Quality_Retrieved_Average_Sigma = "3.255918" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_7\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_7\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_7\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_7\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_7\:Good_Quality = "22" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_7\:Good_Quality_Retrieved = "18" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_7\:Good_Quality_Retrieved_Average_Sigma = "0.561522" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_7\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_7\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_7\:Good_Quality_Failed_Poor_Fit = "4" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_7\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_7\:Good_Quality_Failed_Maxiter = "2" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_7\:Good_Quality_Failed_OOLUT = "1" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_7\:Poor_Quality = "17" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_7\:Poor_Quality_Retrieved = "7" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_7\:Poor_Quality_Retrieved_Average_Sigma = "1.677722" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_8\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_8\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_8\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_8\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_8\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_8\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_8\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_8\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_8\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_8\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_8\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_8\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_8\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_8\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_8\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_8\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_9\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_9\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_9\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_9\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_9\:Good_Quality = "273" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_9\:Good_Quality_Retrieved = "160" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_9\:Good_Quality_Retrieved_Average_Sigma = "2.599082" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_9\:Good_Quality_Failed_Outside_Valid_Range = "33" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_9\:Good_Quality_Failed_Sigma_Too_High = "65" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_9\:Good_Quality_Failed_Poor_Fit = "85" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_9\:Good_Quality_Failed_Marquardt = "13" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_9\:Good_Quality_Failed_Maxiter = "32" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_9\:Good_Quality_Failed_OOLUT = "85" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_9\:Poor_Quality = "288" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_9\:Poor_Quality_Retrieved = "240" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_9\:Poor_Quality_Retrieved_Average_Sigma = "3.081223" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_10\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_10\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_10\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_10\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_10\:Good_Quality = "8069" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_10\:Good_Quality_Retrieved = "5269" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_10\:Good_Quality_Retrieved_Average_Sigma = "2.785885" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_10\:Good_Quality_Failed_Outside_Valid_Range = "379" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_10\:Good_Quality_Failed_Sigma_Too_High = "1082" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_10\:Good_Quality_Failed_Poor_Fit = "2346" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_10\:Good_Quality_Failed_Marquardt = "139" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_10\:Good_Quality_Failed_Maxiter = "195" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_10\:Good_Quality_Failed_OOLUT = "1200" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_10\:Poor_Quality = "1600" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_10\:Poor_Quality_Retrieved = "1075" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_10\:Poor_Quality_Retrieved_Average_Sigma = "3.307963" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_11\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_11\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_11\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_11\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_11\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_11\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_11\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_11\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_11\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_11\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_11\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_11\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_11\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_11\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_11\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_11\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_12\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_12\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_12\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_12\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_12\:Good_Quality = "7009" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_12\:Good_Quality_Retrieved = "5885" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_12\:Good_Quality_Retrieved_Average_Sigma = "1.320947" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_12\:Good_Quality_Failed_Outside_Valid_Range = "4" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_12\:Good_Quality_Failed_Sigma_Too_High = "14" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_12\:Good_Quality_Failed_Poor_Fit = "1027" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_12\:Good_Quality_Failed_Marquardt = "48" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_12\:Good_Quality_Failed_Maxiter = "83" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_12\:Good_Quality_Failed_OOLUT = "38" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_12\:Poor_Quality = "1990" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_12\:Poor_Quality_Retrieved = "1563" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_12\:Poor_Quality_Retrieved_Average_Sigma = "2.000069" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_13\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_13\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_13\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_13\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_13\:Good_Quality = "15933" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_13\:Good_Quality_Retrieved = "13481" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_13\:Good_Quality_Retrieved_Average_Sigma = "1.377319" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_13\:Good_Quality_Failed_Outside_Valid_Range = "22" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_13\:Good_Quality_Failed_Sigma_Too_High = "43" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_13\:Good_Quality_Failed_Poor_Fit = "2414" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_13\:Good_Quality_Failed_Marquardt = "5" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_13\:Good_Quality_Failed_Maxiter = "30" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_13\:Good_Quality_Failed_OOLUT = "72" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_13\:Poor_Quality = "3587" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_13\:Poor_Quality_Retrieved = "2944" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_13\:Poor_Quality_Retrieved_Average_Sigma = "2.700215" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_14\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_14\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_14\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_14\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_14\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_14\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_14\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_14\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_14\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_14\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_14\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_14\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_14\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_14\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_14\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_14\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_15\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_15\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_15\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_15\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_15\:Good_Quality = "4315" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_15\:Good_Quality_Retrieved = "2924" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_15\:Good_Quality_Retrieved_Average_Sigma = "0.768287" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_15\:Good_Quality_Failed_Outside_Valid_Range = "18" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_15\:Good_Quality_Failed_Sigma_Too_High = "16" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_15\:Good_Quality_Failed_Poor_Fit = "1107" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_15\:Good_Quality_Failed_Marquardt = "14" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_15\:Good_Quality_Failed_Maxiter = "410" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_15\:Good_Quality_Failed_OOLUT = "52" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_15\:Poor_Quality = "693" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_15\:Poor_Quality_Retrieved = "426" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_15\:Poor_Quality_Retrieved_Average_Sigma = "1.355604" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_16\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_16\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_16\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_16\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_16\:Good_Quality = "13204" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_16\:Good_Quality_Retrieved = "10058" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_16\:Good_Quality_Retrieved_Average_Sigma = "0.878298" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_16\:Good_Quality_Failed_Outside_Valid_Range = "2" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_16\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_16\:Good_Quality_Failed_Poor_Fit = "3142" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_16\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_16\:Good_Quality_Failed_Maxiter = "29" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_16\:Good_Quality_Failed_OOLUT = "60" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_16\:Poor_Quality = "1291" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_16\:Poor_Quality_Retrieved = "989" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_16\:Poor_Quality_Retrieved_Average_Sigma = "1.659203" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_17\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_17\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_17\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_17\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_17\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_17\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_17\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_17\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_17\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_17\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_17\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_17\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_17\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_17\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_17\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_17\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_18\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_18\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_18\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_18\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_18\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_18\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_18\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_18\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_18\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_18\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_18\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_18\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_18\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_18\:Poor_Quality = "12" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_18\:Poor_Quality_Retrieved = "5" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_18\:Poor_Quality_Retrieved_Average_Sigma = "4.724520" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_19\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_19\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_19\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_19\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_19\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_19\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_19\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_19\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_19\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_19\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_19\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_19\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_19\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_19\:Poor_Quality = "7" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_19\:Poor_Quality_Retrieved = "2" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_19\:Poor_Quality_Retrieved_Average_Sigma = "3.689911" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_20\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_20\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_20\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_20\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_20\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_20\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_20\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_20\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_20\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_20\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_20\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_20\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_20\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_20\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_20\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_20\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_21\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_21\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_21\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_21\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_21\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_21\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_21\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_21\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_21\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_21\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_21\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_21\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_21\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_21\:Poor_Quality = "45" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_21\:Poor_Quality_Retrieved = "37" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_21\:Poor_Quality_Retrieved_Average_Sigma = "3.072677" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_22\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_22\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_22\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_22\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_22\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_22\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_22\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_22\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_22\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_22\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_22\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_22\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_22\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_22\:Poor_Quality = "136" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_22\:Poor_Quality_Retrieved = "92" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_22\:Poor_Quality_Retrieved_Average_Sigma = "3.238413" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_23\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_23\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_23\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_23\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_23\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_23\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_23\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_23\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_23\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_23\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_23\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_23\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_23\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_23\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_23\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_23\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_24\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_24\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_24\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_24\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_24\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_24\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_24\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_24\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_24\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_24\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_24\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_24\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_24\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_24\:Poor_Quality = "92" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_24\:Poor_Quality_Retrieved = "72" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_24\:Poor_Quality_Retrieved_Average_Sigma = "1.981403" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_25\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_25\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_25\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_25\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_25\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_25\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_25\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_25\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_25\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_25\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_25\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_25\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_25\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_25\:Poor_Quality = "161" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_25\:Poor_Quality_Retrieved = "133" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_25\:Poor_Quality_Retrieved_Average_Sigma = "2.019211" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_26\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_26\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_26\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_26\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_26\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_26\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_26\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_26\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_26\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_26\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_26\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_26\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_26\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_26\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_26\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_26\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:SIQ\:Grid_Point_Type = "Sea_Ice" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:SIQ\:SSS_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:SIQ\:SST_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:SIQ\:WS_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:SIQ\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:SIQ\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:SIQ\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:SIQ\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:SIQ\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:SIQ\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:SIQ\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:SIQ\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:SIQ\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:SIQ\:Poor_Quality = "41" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:SIQ\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:SIQ\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:Retrieval_Scheme = "2" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:Land_Rejected = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:Too_Close_To_Land_Rejected = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:Ice_Rejected = "9107" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:Missing_ECMWF_Rejected = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:Too_Few_Measurements_Rejected = "14105" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:Good_Quality_Grid_Points = "49030" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:Poor_Quality_Grid_Points = "10594" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:SQ\:Grid_Point_Type = "Sea" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:SQ\:SSS_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:SQ\:SST_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:SQ\:WS_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:SQ\:Good_Quality = "42416" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:SQ\:Good_Quality_Retrieved = "32650" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:SQ\:Good_Quality_Retrieved_Average_Sigma = "1.309669" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:SQ\:Good_Quality_Failed_Outside_Valid_Range = "126" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:SQ\:Good_Quality_Failed_Sigma_Too_High = "467" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:SQ\:Good_Quality_Failed_Poor_Fit = "9129" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:SQ\:Good_Quality_Failed_Marquardt = "66" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:SQ\:Good_Quality_Failed_Maxiter = "638" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:SQ\:Good_Quality_Failed_OOLUT = "573" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:SQ\:Poor_Quality = "7258" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:SQ\:Poor_Quality_Retrieved = "4970" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:SQ\:Poor_Quality_Retrieved_Average_Sigma = "2.602561" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:NCQ\:Grid_Point_Type = "Near_Coast" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:NCQ\:SSS_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:NCQ\:SST_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:NCQ\:WS_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:NCQ\:Good_Quality = "6614" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:NCQ\:Good_Quality_Retrieved = "3196" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:NCQ\:Good_Quality_Retrieved_Average_Sigma = "2.316276" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:NCQ\:Good_Quality_Failed_Outside_Valid_Range = "354" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:NCQ\:Good_Quality_Failed_Sigma_Too_High = "863" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:NCQ\:Good_Quality_Failed_Poor_Fit = "3116" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:NCQ\:Good_Quality_Failed_Marquardt = "226" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:NCQ\:Good_Quality_Failed_Maxiter = "331" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:NCQ\:Good_Quality_Failed_OOLUT = "1302" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:NCQ\:Poor_Quality = "3336" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:NCQ\:Poor_Quality_Retrieved = "2146" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:NCQ\:Poor_Quality_Retrieved_Average_Sigma = "2.596146" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_0\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_0\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_0\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_0\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_0\:Good_Quality = "40" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_0\:Good_Quality_Retrieved = "10" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_0\:Good_Quality_Retrieved_Average_Sigma = "2.410896" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_0\:Good_Quality_Failed_Outside_Valid_Range = "11" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_0\:Good_Quality_Failed_Sigma_Too_High = "13" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_0\:Good_Quality_Failed_Poor_Fit = "29" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_0\:Good_Quality_Failed_Marquardt = "8" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_0\:Good_Quality_Failed_Maxiter = "3" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_0\:Good_Quality_Failed_OOLUT = "17" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_0\:Poor_Quality = "11" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_0\:Poor_Quality_Retrieved = "5" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_0\:Poor_Quality_Retrieved_Average_Sigma = "4.593025" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_1\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_1\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_1\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_1\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_1\:Good_Quality = "32" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_1\:Good_Quality_Retrieved = "23" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_1\:Good_Quality_Retrieved_Average_Sigma = "2.439510" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_1\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_1\:Good_Quality_Failed_Sigma_Too_High = "3" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_1\:Good_Quality_Failed_Poor_Fit = "9" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_1\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_1\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_1\:Good_Quality_Failed_OOLUT = "6" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_1\:Poor_Quality = "185" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_1\:Poor_Quality_Retrieved = "8" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_1\:Poor_Quality_Retrieved_Average_Sigma = "4.803418" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_2\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_2\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_2\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_2\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_2\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_2\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_2\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_2\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_2\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_2\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_2\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_2\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_2\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_2\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_2\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_2\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_3\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_3\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_3\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_3\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_3\:Good_Quality = "6" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_3\:Good_Quality_Retrieved = "6" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_3\:Good_Quality_Retrieved_Average_Sigma = "1.840680" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_3\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_3\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_3\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_3\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_3\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_3\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_3\:Poor_Quality = "92" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_3\:Poor_Quality_Retrieved = "47" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_3\:Poor_Quality_Retrieved_Average_Sigma = "4.075317" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_4\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_4\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_4\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_4\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_4\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_4\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_4\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_4\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_4\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_4\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_4\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_4\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_4\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_4\:Poor_Quality = "371" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_4\:Poor_Quality_Retrieved = "129" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_4\:Poor_Quality_Retrieved_Average_Sigma = "4.287936" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_5\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_5\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_5\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_5\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_5\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_5\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_5\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_5\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_5\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_5\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_5\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_5\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_5\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_5\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_5\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_5\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_6\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_6\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_6\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_6\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_6\:Good_Quality = "127" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_6\:Good_Quality_Retrieved = "28" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_6\:Good_Quality_Retrieved_Average_Sigma = "0.560374" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_6\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_6\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_6\:Good_Quality_Failed_Poor_Fit = "94" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_6\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_6\:Good_Quality_Failed_Maxiter = "28" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_6\:Good_Quality_Failed_OOLUT = "23" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_6\:Poor_Quality = "16" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_6\:Poor_Quality_Retrieved = "1" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_6\:Poor_Quality_Retrieved_Average_Sigma = "1.426370" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_7\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_7\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_7\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_7\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_7\:Good_Quality = "22" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_7\:Good_Quality_Retrieved = "16" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_7\:Good_Quality_Retrieved_Average_Sigma = "0.547665" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_7\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_7\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_7\:Good_Quality_Failed_Poor_Fit = "6" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_7\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_7\:Good_Quality_Failed_Maxiter = "2" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_7\:Good_Quality_Failed_OOLUT = "1" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_7\:Poor_Quality = "17" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_7\:Poor_Quality_Retrieved = "7" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_7\:Poor_Quality_Retrieved_Average_Sigma = "1.832616" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_8\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_8\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_8\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_8\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_8\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_8\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_8\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_8\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_8\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_8\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_8\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_8\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_8\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_8\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_8\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_8\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_9\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_9\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_9\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_9\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_9\:Good_Quality = "273" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_9\:Good_Quality_Retrieved = "155" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_9\:Good_Quality_Retrieved_Average_Sigma = "2.577458" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_9\:Good_Quality_Failed_Outside_Valid_Range = "35" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_9\:Good_Quality_Failed_Sigma_Too_High = "68" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_9\:Good_Quality_Failed_Poor_Fit = "86" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_9\:Good_Quality_Failed_Marquardt = "14" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_9\:Good_Quality_Failed_Maxiter = "34" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_9\:Good_Quality_Failed_OOLUT = "89" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_9\:Poor_Quality = "288" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_9\:Poor_Quality_Retrieved = "244" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_9\:Poor_Quality_Retrieved_Average_Sigma = "3.173979" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_10\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_10\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_10\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_10\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_10\:Good_Quality = "8069" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_10\:Good_Quality_Retrieved = "5009" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_10\:Good_Quality_Retrieved_Average_Sigma = "2.802226" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_10\:Good_Quality_Failed_Outside_Valid_Range = "381" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_10\:Good_Quality_Failed_Sigma_Too_High = "1149" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_10\:Good_Quality_Failed_Poor_Fit = "2608" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_10\:Good_Quality_Failed_Marquardt = "146" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_10\:Good_Quality_Failed_Maxiter = "192" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_10\:Good_Quality_Failed_OOLUT = "1331" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_10\:Poor_Quality = "1600" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_10\:Poor_Quality_Retrieved = "1041" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_10\:Poor_Quality_Retrieved_Average_Sigma = "3.312484" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_11\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_11\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_11\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_11\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_11\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_11\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_11\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_11\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_11\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_11\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_11\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_11\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_11\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_11\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_11\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_11\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_12\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_12\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_12\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_12\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_12\:Good_Quality = "7009" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_12\:Good_Quality_Retrieved = "5553" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_12\:Good_Quality_Retrieved_Average_Sigma = "1.349544" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_12\:Good_Quality_Failed_Outside_Valid_Range = "8" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_12\:Good_Quality_Failed_Sigma_Too_High = "19" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_12\:Good_Quality_Failed_Poor_Fit = "1358" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_12\:Good_Quality_Failed_Marquardt = "70" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_12\:Good_Quality_Failed_Maxiter = "126" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_12\:Good_Quality_Failed_OOLUT = "68" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_12\:Poor_Quality = "1990" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_12\:Poor_Quality_Retrieved = "1438" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_12\:Poor_Quality_Retrieved_Average_Sigma = "2.169792" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_13\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_13\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_13\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_13\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_13\:Good_Quality = "15933" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_13\:Good_Quality_Retrieved = "12618" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_13\:Good_Quality_Retrieved_Average_Sigma = "1.389448" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_13\:Good_Quality_Failed_Outside_Valid_Range = "16" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_13\:Good_Quality_Failed_Sigma_Too_High = "48" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_13\:Good_Quality_Failed_Poor_Fit = "3254" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_13\:Good_Quality_Failed_Marquardt = "11" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_13\:Good_Quality_Failed_Maxiter = "79" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_13\:Good_Quality_Failed_OOLUT = "214" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_13\:Poor_Quality = "3587" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_13\:Poor_Quality_Retrieved = "2533" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_13\:Poor_Quality_Retrieved_Average_Sigma = "2.911479" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_14\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_14\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_14\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_14\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_14\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_14\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_14\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_14\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_14\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_14\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_14\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_14\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_14\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_14\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_14\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_14\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_15\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_15\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_15\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_15\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_15\:Good_Quality = "4315" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_15\:Good_Quality_Retrieved = "2837" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_15\:Good_Quality_Retrieved_Average_Sigma = "0.767496" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_15\:Good_Quality_Failed_Outside_Valid_Range = "29" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_15\:Good_Quality_Failed_Sigma_Too_High = "30" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_15\:Good_Quality_Failed_Poor_Fit = "1196" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_15\:Good_Quality_Failed_Marquardt = "43" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_15\:Good_Quality_Failed_Maxiter = "474" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_15\:Good_Quality_Failed_OOLUT = "67" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_15\:Poor_Quality = "693" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_15\:Poor_Quality_Retrieved = "404" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_15\:Poor_Quality_Retrieved_Average_Sigma = "1.257553" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_16\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_16\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_16\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_16\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_16\:Good_Quality = "13204" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_16\:Good_Quality_Retrieved = "9591" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_16\:Good_Quality_Retrieved_Average_Sigma = "0.876707" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_16\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_16\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_16\:Good_Quality_Failed_Poor_Fit = "3605" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_16\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_16\:Good_Quality_Failed_Maxiter = "31" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_16\:Good_Quality_Failed_OOLUT = "59" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_16\:Poor_Quality = "1291" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_16\:Poor_Quality_Retrieved = "907" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_16\:Poor_Quality_Retrieved_Average_Sigma = "1.710565" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_17\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_17\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_17\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_17\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_17\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_17\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_17\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_17\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_17\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_17\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_17\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_17\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_17\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_17\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_17\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_17\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_18\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_18\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_18\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_18\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_18\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_18\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_18\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_18\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_18\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_18\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_18\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_18\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_18\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_18\:Poor_Quality = "12" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_18\:Poor_Quality_Retrieved = "5" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_18\:Poor_Quality_Retrieved_Average_Sigma = "4.715192" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_19\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_19\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_19\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_19\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_19\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_19\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_19\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_19\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_19\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_19\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_19\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_19\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_19\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_19\:Poor_Quality = "7" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_19\:Poor_Quality_Retrieved = "2" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_19\:Poor_Quality_Retrieved_Average_Sigma = "3.695637" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_20\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_20\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_20\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_20\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_20\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_20\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_20\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_20\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_20\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_20\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_20\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_20\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_20\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_20\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_20\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_20\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_21\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_21\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_21\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_21\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_21\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_21\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_21\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_21\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_21\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_21\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_21\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_21\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_21\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_21\:Poor_Quality = "45" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_21\:Poor_Quality_Retrieved = "34" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_21\:Poor_Quality_Retrieved_Average_Sigma = "3.077266" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_22\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_22\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_22\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_22\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_22\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_22\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_22\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_22\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_22\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_22\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_22\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_22\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_22\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_22\:Poor_Quality = "136" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_22\:Poor_Quality_Retrieved = "104" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_22\:Poor_Quality_Retrieved_Average_Sigma = "3.421102" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_23\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_23\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_23\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_23\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_23\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_23\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_23\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_23\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_23\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_23\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_23\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_23\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_23\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_23\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_23\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_23\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_24\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_24\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_24\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_24\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_24\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_24\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_24\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_24\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_24\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_24\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_24\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_24\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_24\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_24\:Poor_Quality = "92" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_24\:Poor_Quality_Retrieved = "74" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_24\:Poor_Quality_Retrieved_Average_Sigma = "2.013027" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_25\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_25\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_25\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_25\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_25\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_25\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_25\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_25\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_25\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_25\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_25\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_25\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_25\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_25\:Poor_Quality = "161" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_25\:Poor_Quality_Retrieved = "133" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_25\:Poor_Quality_Retrieved_Average_Sigma = "2.016223" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_26\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_26\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_26\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_26\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_26\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_26\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_26\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_26\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_26\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_26\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_26\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_26\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_26\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_26\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_26\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_26\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:SIQ\:Grid_Point_Type = "Sea_Ice" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:SIQ\:SSS_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:SIQ\:SST_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:SIQ\:WS_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:SIQ\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:SIQ\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:SIQ\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:SIQ\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:SIQ\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:SIQ\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:SIQ\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:SIQ\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:SIQ\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:SIQ\:Poor_Quality = "41" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:SIQ\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:SIQ\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:Retrieval_Scheme = "3" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:Land_Rejected = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:Too_Close_To_Land_Rejected = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:Ice_Rejected = "9107" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:Missing_ECMWF_Rejected = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:Too_Few_Measurements_Rejected = "14105" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:Good_Quality_Grid_Points = "49030" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:Poor_Quality_Grid_Points = "10594" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:SQ\:Grid_Point_Type = "Sea" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:SQ\:SSS_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:SQ\:SST_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:SQ\:WS_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:SQ\:Good_Quality = "42416" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:SQ\:Good_Quality_Retrieved = "33881" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:SQ\:Good_Quality_Retrieved_Average_Sigma = "1.300973" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:SQ\:Good_Quality_Failed_Outside_Valid_Range = "138" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:SQ\:Good_Quality_Failed_Sigma_Too_High = "456" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:SQ\:Good_Quality_Failed_Poor_Fit = "7974" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:SQ\:Good_Quality_Failed_Marquardt = "50" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:SQ\:Good_Quality_Failed_Maxiter = "489" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:SQ\:Good_Quality_Failed_OOLUT = "549" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:SQ\:Poor_Quality = "7258" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:SQ\:Poor_Quality_Retrieved = "5481" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:SQ\:Poor_Quality_Retrieved_Average_Sigma = "2.500925" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:NCQ\:Grid_Point_Type = "Near_Coast" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:NCQ\:SSS_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:NCQ\:SST_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:NCQ\:WS_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:NCQ\:Good_Quality = "6614" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:NCQ\:Good_Quality_Retrieved = "3994" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:NCQ\:Good_Quality_Retrieved_Average_Sigma = "2.145041" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:NCQ\:Good_Quality_Failed_Outside_Valid_Range = "331" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:NCQ\:Good_Quality_Failed_Sigma_Too_High = "780" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:NCQ\:Good_Quality_Failed_Poor_Fit = "2270" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:NCQ\:Good_Quality_Failed_Marquardt = "175" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:NCQ\:Good_Quality_Failed_Maxiter = "307" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:NCQ\:Good_Quality_Failed_OOLUT = "993" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:NCQ\:Poor_Quality = "3336" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:NCQ\:Poor_Quality_Retrieved = "2402" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:NCQ\:Poor_Quality_Retrieved_Average_Sigma = "2.491391" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_0\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_0\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_0\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_0\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_0\:Good_Quality = "40" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_0\:Good_Quality_Retrieved = "13" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_0\:Good_Quality_Retrieved_Average_Sigma = "2.271775" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_0\:Good_Quality_Failed_Outside_Valid_Range = "11" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_0\:Good_Quality_Failed_Sigma_Too_High = "13" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_0\:Good_Quality_Failed_Poor_Fit = "26" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_0\:Good_Quality_Failed_Marquardt = "6" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_0\:Good_Quality_Failed_Maxiter = "6" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_0\:Good_Quality_Failed_OOLUT = "14" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_0\:Poor_Quality = "11" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_0\:Poor_Quality_Retrieved = "6" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_0\:Poor_Quality_Retrieved_Average_Sigma = "4.644665" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_1\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_1\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_1\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_1\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_1\:Good_Quality = "32" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_1\:Good_Quality_Retrieved = "25" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_1\:Good_Quality_Retrieved_Average_Sigma = "2.331885" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_1\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_1\:Good_Quality_Failed_Sigma_Too_High = "3" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_1\:Good_Quality_Failed_Poor_Fit = "6" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_1\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_1\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_1\:Good_Quality_Failed_OOLUT = "4" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_1\:Poor_Quality = "185" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_1\:Poor_Quality_Retrieved = "8" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_1\:Poor_Quality_Retrieved_Average_Sigma = "4.768177" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_2\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_2\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_2\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_2\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_2\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_2\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_2\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_2\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_2\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_2\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_2\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_2\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_2\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_2\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_2\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_2\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_3\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_3\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_3\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_3\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_3\:Good_Quality = "6" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_3\:Good_Quality_Retrieved = "6" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_3\:Good_Quality_Retrieved_Average_Sigma = "1.849856" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_3\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_3\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_3\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_3\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_3\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_3\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_3\:Poor_Quality = "92" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_3\:Poor_Quality_Retrieved = "61" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_3\:Poor_Quality_Retrieved_Average_Sigma = "3.938132" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_4\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_4\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_4\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_4\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_4\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_4\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_4\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_4\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_4\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_4\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_4\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_4\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_4\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_4\:Poor_Quality = "371" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_4\:Poor_Quality_Retrieved = "214" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_4\:Poor_Quality_Retrieved_Average_Sigma = "4.211347" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_5\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_5\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_5\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_5\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_5\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_5\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_5\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_5\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_5\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_5\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_5\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_5\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_5\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_5\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_5\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_5\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_6\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_6\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_6\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_6\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_6\:Good_Quality = "127" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_6\:Good_Quality_Retrieved = "36" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_6\:Good_Quality_Retrieved_Average_Sigma = "0.556612" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_6\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_6\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_6\:Good_Quality_Failed_Poor_Fit = "87" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_6\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_6\:Good_Quality_Failed_Maxiter = "9" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_6\:Good_Quality_Failed_OOLUT = "16" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_6\:Poor_Quality = "16" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_6\:Poor_Quality_Retrieved = "9" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_6\:Poor_Quality_Retrieved_Average_Sigma = "3.255918" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_7\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_7\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_7\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_7\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_7\:Good_Quality = "22" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_7\:Good_Quality_Retrieved = "18" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_7\:Good_Quality_Retrieved_Average_Sigma = "0.561522" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_7\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_7\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_7\:Good_Quality_Failed_Poor_Fit = "4" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_7\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_7\:Good_Quality_Failed_Maxiter = "2" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_7\:Good_Quality_Failed_OOLUT = "1" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_7\:Poor_Quality = "17" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_7\:Poor_Quality_Retrieved = "7" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_7\:Poor_Quality_Retrieved_Average_Sigma = "1.677722" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_8\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_8\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_8\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_8\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_8\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_8\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_8\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_8\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_8\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_8\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_8\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_8\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_8\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_8\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_8\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_8\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_9\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_9\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_9\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_9\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_9\:Good_Quality = "273" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_9\:Good_Quality_Retrieved = "160" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_9\:Good_Quality_Retrieved_Average_Sigma = "2.599082" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_9\:Good_Quality_Failed_Outside_Valid_Range = "33" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_9\:Good_Quality_Failed_Sigma_Too_High = "65" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_9\:Good_Quality_Failed_Poor_Fit = "85" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_9\:Good_Quality_Failed_Marquardt = "13" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_9\:Good_Quality_Failed_Maxiter = "32" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_9\:Good_Quality_Failed_OOLUT = "85" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_9\:Poor_Quality = "288" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_9\:Poor_Quality_Retrieved = "240" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_9\:Poor_Quality_Retrieved_Average_Sigma = "3.081223" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_10\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_10\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_10\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_10\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_10\:Good_Quality = "8069" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_10\:Good_Quality_Retrieved = "5269" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_10\:Good_Quality_Retrieved_Average_Sigma = "2.785885" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_10\:Good_Quality_Failed_Outside_Valid_Range = "379" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_10\:Good_Quality_Failed_Sigma_Too_High = "1082" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_10\:Good_Quality_Failed_Poor_Fit = "2346" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_10\:Good_Quality_Failed_Marquardt = "139" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_10\:Good_Quality_Failed_Maxiter = "195" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_10\:Good_Quality_Failed_OOLUT = "1200" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_10\:Poor_Quality = "1600" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_10\:Poor_Quality_Retrieved = "1075" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_10\:Poor_Quality_Retrieved_Average_Sigma = "3.307963" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_11\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_11\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_11\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_11\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_11\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_11\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_11\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_11\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_11\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_11\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_11\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_11\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_11\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_11\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_11\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_11\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_12\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_12\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_12\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_12\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_12\:Good_Quality = "7009" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_12\:Good_Quality_Retrieved = "5885" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_12\:Good_Quality_Retrieved_Average_Sigma = "1.320947" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_12\:Good_Quality_Failed_Outside_Valid_Range = "4" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_12\:Good_Quality_Failed_Sigma_Too_High = "14" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_12\:Good_Quality_Failed_Poor_Fit = "1027" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_12\:Good_Quality_Failed_Marquardt = "48" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_12\:Good_Quality_Failed_Maxiter = "83" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_12\:Good_Quality_Failed_OOLUT = "38" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_12\:Poor_Quality = "1990" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_12\:Poor_Quality_Retrieved = "1563" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_12\:Poor_Quality_Retrieved_Average_Sigma = "2.000069" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_13\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_13\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_13\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_13\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_13\:Good_Quality = "15933" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_13\:Good_Quality_Retrieved = "13481" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_13\:Good_Quality_Retrieved_Average_Sigma = "1.377319" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_13\:Good_Quality_Failed_Outside_Valid_Range = "22" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_13\:Good_Quality_Failed_Sigma_Too_High = "43" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_13\:Good_Quality_Failed_Poor_Fit = "2414" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_13\:Good_Quality_Failed_Marquardt = "5" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_13\:Good_Quality_Failed_Maxiter = "30" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_13\:Good_Quality_Failed_OOLUT = "72" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_13\:Poor_Quality = "3587" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_13\:Poor_Quality_Retrieved = "2944" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_13\:Poor_Quality_Retrieved_Average_Sigma = "2.700215" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_14\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_14\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_14\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_14\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_14\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_14\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_14\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_14\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_14\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_14\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_14\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_14\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_14\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_14\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_14\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_14\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_15\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_15\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_15\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_15\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_15\:Good_Quality = "4315" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_15\:Good_Quality_Retrieved = "2924" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_15\:Good_Quality_Retrieved_Average_Sigma = "0.768287" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_15\:Good_Quality_Failed_Outside_Valid_Range = "18" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_15\:Good_Quality_Failed_Sigma_Too_High = "16" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_15\:Good_Quality_Failed_Poor_Fit = "1107" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_15\:Good_Quality_Failed_Marquardt = "14" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_15\:Good_Quality_Failed_Maxiter = "410" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_15\:Good_Quality_Failed_OOLUT = "52" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_15\:Poor_Quality = "693" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_15\:Poor_Quality_Retrieved = "426" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_15\:Poor_Quality_Retrieved_Average_Sigma = "1.355604" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_16\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_16\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_16\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_16\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_16\:Good_Quality = "13204" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_16\:Good_Quality_Retrieved = "10058" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_16\:Good_Quality_Retrieved_Average_Sigma = "0.878298" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_16\:Good_Quality_Failed_Outside_Valid_Range = "2" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_16\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_16\:Good_Quality_Failed_Poor_Fit = "3142" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_16\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_16\:Good_Quality_Failed_Maxiter = "29" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_16\:Good_Quality_Failed_OOLUT = "60" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_16\:Poor_Quality = "1291" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_16\:Poor_Quality_Retrieved = "989" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_16\:Poor_Quality_Retrieved_Average_Sigma = "1.659203" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_17\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_17\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_17\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_17\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_17\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_17\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_17\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_17\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_17\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_17\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_17\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_17\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_17\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_17\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_17\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_17\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_18\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_18\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_18\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_18\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_18\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_18\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_18\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_18\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_18\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_18\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_18\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_18\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_18\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_18\:Poor_Quality = "12" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_18\:Poor_Quality_Retrieved = "5" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_18\:Poor_Quality_Retrieved_Average_Sigma = "4.724520" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_19\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_19\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_19\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_19\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_19\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_19\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_19\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_19\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_19\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_19\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_19\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_19\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_19\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_19\:Poor_Quality = "7" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_19\:Poor_Quality_Retrieved = "2" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_19\:Poor_Quality_Retrieved_Average_Sigma = "3.689911" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_20\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_20\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_20\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_20\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_20\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_20\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_20\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_20\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_20\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_20\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_20\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_20\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_20\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_20\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_20\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_20\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_21\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_21\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_21\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_21\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_21\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_21\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_21\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_21\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_21\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_21\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_21\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_21\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_21\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_21\:Poor_Quality = "45" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_21\:Poor_Quality_Retrieved = "37" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_21\:Poor_Quality_Retrieved_Average_Sigma = "3.072677" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_22\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_22\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_22\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_22\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_22\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_22\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_22\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_22\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_22\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_22\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_22\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_22\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_22\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_22\:Poor_Quality = "136" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_22\:Poor_Quality_Retrieved = "92" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_22\:Poor_Quality_Retrieved_Average_Sigma = "3.238413" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_23\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_23\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_23\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_23\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_23\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_23\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_23\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_23\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_23\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_23\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_23\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_23\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_23\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_23\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_23\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_23\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_24\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_24\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_24\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_24\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_24\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_24\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_24\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_24\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_24\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_24\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_24\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_24\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_24\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_24\:Poor_Quality = "92" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_24\:Poor_Quality_Retrieved = "72" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_24\:Poor_Quality_Retrieved_Average_Sigma = "1.981403" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_25\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_25\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_25\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_25\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_25\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_25\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_25\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_25\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_25\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_25\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_25\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_25\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_25\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_25\:Poor_Quality = "161" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_25\:Poor_Quality_Retrieved = "133" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_25\:Poor_Quality_Retrieved_Average_Sigma = "2.019211" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_26\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_26\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_26\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_26\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_26\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_26\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_26\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_26\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_26\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_26\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_26\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_26\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_26\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_26\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_26\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_26\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:SIQ\:Grid_Point_Type = "Sea_Ice" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:SIQ\:SSS_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:SIQ\:SST_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:SIQ\:WS_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:SIQ\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:SIQ\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:SIQ\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:SIQ\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:SIQ\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:SIQ\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:SIQ\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:SIQ\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:SIQ\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:SIQ\:Poor_Quality = "41" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:SIQ\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:SIQ\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:Retrieval_Scheme = "4" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:Land_Rejected = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:Too_Close_To_Land_Rejected = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:Ice_Rejected = "9107" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:Missing_ECMWF_Rejected = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:Too_Few_Measurements_Rejected = "14105" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:Good_Quality_Grid_Points = "49030" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:Poor_Quality_Grid_Points = "10594" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:SQ\:Grid_Point_Type = "Sea" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:SQ\:SSS_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:SQ\:SST_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:SQ\:WS_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:SQ\:Good_Quality = "42416" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:SQ\:Good_Quality_Retrieved = "38092" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:SQ\:Good_Quality_Retrieved_Average_Sigma = "0.777640" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:SQ\:Good_Quality_Failed_Outside_Valid_Range = "725" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:SQ\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:SQ\:Good_Quality_Failed_Poor_Fit = "3680" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:SQ\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:SQ\:Good_Quality_Failed_Maxiter = "5" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:SQ\:Good_Quality_Failed_OOLUT = "3670" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:SQ\:Poor_Quality = "7258" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:SQ\:Poor_Quality_Retrieved = "5930" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:SQ\:Poor_Quality_Retrieved_Average_Sigma = "1.312244" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:NCQ\:Grid_Point_Type = "Near_Coast" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:NCQ\:SSS_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:NCQ\:SST_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:NCQ\:WS_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:NCQ\:Good_Quality = "6614" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:NCQ\:Good_Quality_Retrieved = "5275" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:NCQ\:Good_Quality_Retrieved_Average_Sigma = "0.713190" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:NCQ\:Good_Quality_Failed_Outside_Valid_Range = "108" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:NCQ\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:NCQ\:Good_Quality_Failed_Poor_Fit = "1336" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:NCQ\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:NCQ\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:NCQ\:Good_Quality_Failed_OOLUT = "1330" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:NCQ\:Poor_Quality = "3336" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:NCQ\:Poor_Quality_Retrieved = "2822" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:NCQ\:Poor_Quality_Retrieved_Average_Sigma = "1.012104" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_0\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_0\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_0\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_0\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_0\:Good_Quality = "40" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_0\:Good_Quality_Retrieved = "31" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_0\:Good_Quality_Retrieved_Average_Sigma = "0.584082" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_0\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_0\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_0\:Good_Quality_Failed_Poor_Fit = "9" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_0\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_0\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_0\:Good_Quality_Failed_OOLUT = "9" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_0\:Poor_Quality = "11" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_0\:Poor_Quality_Retrieved = "11" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_0\:Poor_Quality_Retrieved_Average_Sigma = "1.497783" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_1\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_1\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_1\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_1\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_1\:Good_Quality = "32" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_1\:Good_Quality_Retrieved = "30" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_1\:Good_Quality_Retrieved_Average_Sigma = "0.623371" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_1\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_1\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_1\:Good_Quality_Failed_Poor_Fit = "2" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_1\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_1\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_1\:Good_Quality_Failed_OOLUT = "2" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_1\:Poor_Quality = "185" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_1\:Poor_Quality_Retrieved = "120" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_1\:Poor_Quality_Retrieved_Average_Sigma = "1.599651" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_2\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_2\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_2\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_2\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_2\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_2\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_2\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_2\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_2\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_2\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_2\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_2\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_2\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_2\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_2\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_2\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_3\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_3\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_3\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_3\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_3\:Good_Quality = "6" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_3\:Good_Quality_Retrieved = "6" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_3\:Good_Quality_Retrieved_Average_Sigma = "0.953346" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_3\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_3\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_3\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_3\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_3\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_3\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_3\:Poor_Quality = "92" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_3\:Poor_Quality_Retrieved = "72" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_3\:Poor_Quality_Retrieved_Average_Sigma = "1.688501" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_4\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_4\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_4\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_4\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_4\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_4\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_4\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_4\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_4\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_4\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_4\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_4\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_4\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_4\:Poor_Quality = "371" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_4\:Poor_Quality_Retrieved = "314" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_4\:Poor_Quality_Retrieved_Average_Sigma = "1.663750" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_5\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_5\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_5\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_5\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_5\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_5\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_5\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_5\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_5\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_5\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_5\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_5\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_5\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_5\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_5\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_5\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_6\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_6\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_6\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_6\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_6\:Good_Quality = "127" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_6\:Good_Quality_Retrieved = "48" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_6\:Good_Quality_Retrieved_Average_Sigma = "0.726662" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_6\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_6\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_6\:Good_Quality_Failed_Poor_Fit = "79" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_6\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_6\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_6\:Good_Quality_Failed_OOLUT = "79" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_6\:Poor_Quality = "16" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_6\:Poor_Quality_Retrieved = "9" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_6\:Poor_Quality_Retrieved_Average_Sigma = "1.440257" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_7\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_7\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_7\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_7\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_7\:Good_Quality = "22" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_7\:Good_Quality_Retrieved = "18" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_7\:Good_Quality_Retrieved_Average_Sigma = "0.760549" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_7\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_7\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_7\:Good_Quality_Failed_Poor_Fit = "4" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_7\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_7\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_7\:Good_Quality_Failed_OOLUT = "4" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_7\:Poor_Quality = "17" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_7\:Poor_Quality_Retrieved = "6" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_7\:Poor_Quality_Retrieved_Average_Sigma = "1.655105" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_8\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_8\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_8\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_8\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_8\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_8\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_8\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_8\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_8\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_8\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_8\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_8\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_8\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_8\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_8\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_8\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_9\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_9\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_9\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_9\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_9\:Good_Quality = "273" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_9\:Good_Quality_Retrieved = "228" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_9\:Good_Quality_Retrieved_Average_Sigma = "0.667519" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_9\:Good_Quality_Failed_Outside_Valid_Range = "1" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_9\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_9\:Good_Quality_Failed_Poor_Fit = "44" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_9\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_9\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_9\:Good_Quality_Failed_OOLUT = "45" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_9\:Poor_Quality = "288" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_9\:Poor_Quality_Retrieved = "249" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_9\:Poor_Quality_Retrieved_Average_Sigma = "1.094154" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_10\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_10\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_10\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_10\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_10\:Good_Quality = "8069" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_10\:Good_Quality_Retrieved = "6840" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_10\:Good_Quality_Retrieved_Average_Sigma = "0.689680" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_10\:Good_Quality_Failed_Outside_Valid_Range = "83" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_10\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_10\:Good_Quality_Failed_Poor_Fit = "1224" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_10\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_10\:Good_Quality_Failed_Maxiter = "5" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_10\:Good_Quality_Failed_OOLUT = "1229" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_10\:Poor_Quality = "1600" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_10\:Poor_Quality_Retrieved = "1347" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_10\:Poor_Quality_Retrieved_Average_Sigma = "1.023891" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_11\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_11\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_11\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_11\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_11\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_11\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_11\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_11\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_11\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_11\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_11\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_11\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_11\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_11\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_11\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_11\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_12\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_12\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_12\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_12\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_12\:Good_Quality = "7009" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_12\:Good_Quality_Retrieved = "6588" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_12\:Good_Quality_Retrieved_Average_Sigma = "0.757073" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_12\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_12\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_12\:Good_Quality_Failed_Poor_Fit = "421" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_12\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_12\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_12\:Good_Quality_Failed_OOLUT = "414" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_12\:Poor_Quality = "1990" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_12\:Poor_Quality_Retrieved = "1804" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_12\:Poor_Quality_Retrieved_Average_Sigma = "0.902115" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_13\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_13\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_13\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_13\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_13\:Good_Quality = "15933" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_13\:Good_Quality_Retrieved = "14872" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_13\:Good_Quality_Retrieved_Average_Sigma = "0.744029" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_13\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_13\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_13\:Good_Quality_Failed_Poor_Fit = "1061" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_13\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_13\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_13\:Good_Quality_Failed_OOLUT = "1017" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_13\:Poor_Quality = "3587" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_13\:Poor_Quality_Retrieved = "3124" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_13\:Poor_Quality_Retrieved_Average_Sigma = "1.219597" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_14\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_14\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_14\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_14\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_14\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_14\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_14\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_14\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_14\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_14\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_14\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_14\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_14\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_14\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_14\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_14\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_15\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_15\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_15\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_15\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_15\:Good_Quality = "4315" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_15\:Good_Quality_Retrieved = "3022" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_15\:Good_Quality_Retrieved_Average_Sigma = "0.822249" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_15\:Good_Quality_Failed_Outside_Valid_Range = "694" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_15\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_15\:Good_Quality_Failed_Poor_Fit = "675" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_15\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_15\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_15\:Good_Quality_Failed_OOLUT = "1096" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_15\:Poor_Quality = "693" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_15\:Poor_Quality_Retrieved = "418" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_15\:Poor_Quality_Retrieved_Average_Sigma = "1.274173" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_16\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_16\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_16\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_16\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_16\:Good_Quality = "13204" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_16\:Good_Quality_Retrieved = "11684" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_16\:Good_Quality_Retrieved_Average_Sigma = "0.846080" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_16\:Good_Quality_Failed_Outside_Valid_Range = "55" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_16\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_16\:Good_Quality_Failed_Poor_Fit = "1497" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_16\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_16\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_16\:Good_Quality_Failed_OOLUT = "1105" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_16\:Poor_Quality = "1291" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_16\:Poor_Quality_Retrieved = "996" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_16\:Poor_Quality_Retrieved_Average_Sigma = "1.601620" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_17\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_17\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_17\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_17\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_17\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_17\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_17\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_17\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_17\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_17\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_17\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_17\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_17\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_17\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_17\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_17\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_18\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_18\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_18\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_18\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_18\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_18\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_18\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_18\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_18\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_18\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_18\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_18\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_18\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_18\:Poor_Quality = "12" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_18\:Poor_Quality_Retrieved = "9" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_18\:Poor_Quality_Retrieved_Average_Sigma = "1.653254" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_19\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_19\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_19\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_19\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_19\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_19\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_19\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_19\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_19\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_19\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_19\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_19\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_19\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_19\:Poor_Quality = "7" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_19\:Poor_Quality_Retrieved = "6" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_19\:Poor_Quality_Retrieved_Average_Sigma = "1.644945" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_20\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_20\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_20\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_20\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_20\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_20\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_20\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_20\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_20\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_20\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_20\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_20\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_20\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_20\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_20\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_20\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_21\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_21\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_21\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_21\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_21\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_21\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_21\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_21\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_21\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_21\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_21\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_21\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_21\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_21\:Poor_Quality = "45" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_21\:Poor_Quality_Retrieved = "41" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_21\:Poor_Quality_Retrieved_Average_Sigma = "1.816824" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_22\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_22\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_22\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_22\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_22\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_22\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_22\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_22\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_22\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_22\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_22\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_22\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_22\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_22\:Poor_Quality = "136" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_22\:Poor_Quality_Retrieved = "102" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_22\:Poor_Quality_Retrieved_Average_Sigma = "1.893596" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_23\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_23\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_23\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_23\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_23\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_23\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_23\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_23\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_23\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_23\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_23\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_23\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_23\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_23\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_23\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_23\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_24\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_24\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_24\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_24\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_24\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_24\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_24\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_24\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_24\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_24\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_24\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_24\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_24\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_24\:Poor_Quality = "92" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_24\:Poor_Quality_Retrieved = "31" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_24\:Poor_Quality_Retrieved_Average_Sigma = "2.030431" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_25\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_25\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_25\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_25\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_25\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_25\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_25\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_25\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_25\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_25\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_25\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_25\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_25\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_25\:Poor_Quality = "161" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_25\:Poor_Quality_Retrieved = "93" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_25\:Poor_Quality_Retrieved_Average_Sigma = "2.045601" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_26\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_26\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_26\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_26\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_26\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_26\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_26\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_26\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_26\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_26\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_26\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_26\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_26\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_26\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_26\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_26\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:SIQ\:Grid_Point_Type = "Sea_Ice" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:SIQ\:SSS_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:SIQ\:SST_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:SIQ\:WS_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:SIQ\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:SIQ\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:SIQ\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:SIQ\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:SIQ\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:SIQ\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:SIQ\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:SIQ\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:SIQ\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:SIQ\:Poor_Quality = "41" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:SIQ\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:SIQ\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_0\:Retrieved_Parameter_0\:name = "SSS" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_0\:Retrieved_Parameter_0\:unit = "Practical Salinity Unit (PSU)" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_0\:Retrieved_Parameter_0\:description = "Surface salinity of the sea at gridpoint" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_0\:Retrieved_Parameter_1\:name = "SST" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_0\:Retrieved_Parameter_1\:unit = "Kelvin" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_0\:Retrieved_Parameter_1\:description = "Surface temperature of the sea at gridpoint" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_0\:Retrieved_Parameter_2\:name = "UN10" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_0\:Retrieved_Parameter_2\:unit = "m.s-1" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_0\:Retrieved_Parameter_2\:description = "U component of neutral wind 10m above surface" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_0\:Retrieved_Parameter_3\:name = "VN10" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_0\:Retrieved_Parameter_3\:unit = "m.s-1" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_0\:Retrieved_Parameter_3\:description = "V component of neutral wind 10m above surface" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_0\:Retrieved_Parameter_4\:name = "tec" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_0\:Retrieved_Parameter_4\:unit = "tecu" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_0\:Retrieved_Parameter_4\:description = "Total Electronic Content of the ionosphere below SMOS" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_0\:Retrieved_Parameter_5\:name = "not used" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_0\:Retrieved_Parameter_5\:unit = "none" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_0\:Retrieved_Parameter_5\:description = "no parameter defined" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_0\:Retrieved_Parameter_6\:name = "not used" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_0\:Retrieved_Parameter_6\:unit = "none" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_0\:Retrieved_Parameter_6\:description = "no parameter defined" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_0\:Retrieved_Parameter_7\:name = "not used" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_0\:Retrieved_Parameter_7\:unit = "none" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_0\:Retrieved_Parameter_7\:description = "no parameter defined" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_0\:Retrieved_Parameter_8\:name = "not used" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_0\:Retrieved_Parameter_8\:unit = "none" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_0\:Retrieved_Parameter_8\:description = "no parameter defined" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_0\:Retrieved_Parameter_9\:name = "not used" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_0\:Retrieved_Parameter_9\:unit = "none" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_0\:Retrieved_Parameter_9\:description = "no parameter defined" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_1\:Retrieved_Parameter_0\:name = "SSS" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_1\:Retrieved_Parameter_0\:unit = "Practical Salinity Unit (PSU)" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_1\:Retrieved_Parameter_0\:description = "Surface salinity of the sea at gridpoint" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_1\:Retrieved_Parameter_1\:name = "SST" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_1\:Retrieved_Parameter_1\:unit = "Kelvin" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_1\:Retrieved_Parameter_1\:description = "Surface temperature of the sea at gridpoint" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_1\:Retrieved_Parameter_2\:name = "UN10" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_1\:Retrieved_Parameter_2\:unit = "m.s-1" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_1\:Retrieved_Parameter_2\:description = "U component of neutral wind 10m above surface" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_1\:Retrieved_Parameter_3\:name = "VN10" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_1\:Retrieved_Parameter_3\:unit = "m.s-1" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_1\:Retrieved_Parameter_3\:description = "V component of neutral wind 10m above surface" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_1\:Retrieved_Parameter_4\:name = "tec" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_1\:Retrieved_Parameter_4\:unit = "tecu" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_1\:Retrieved_Parameter_4\:description = "Total Electronic Content of the ionosphere below SMOS" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_1\:Retrieved_Parameter_5\:name = "not used" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_1\:Retrieved_Parameter_5\:unit = "none" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_1\:Retrieved_Parameter_5\:description = "no parameter defined" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_1\:Retrieved_Parameter_6\:name = "not used" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_1\:Retrieved_Parameter_6\:unit = "none" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_1\:Retrieved_Parameter_6\:description = "no parameter defined" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_1\:Retrieved_Parameter_7\:name = "not used" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_1\:Retrieved_Parameter_7\:unit = "none" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_1\:Retrieved_Parameter_7\:description = "no parameter defined" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_1\:Retrieved_Parameter_8\:name = "not used" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_1\:Retrieved_Parameter_8\:unit = "none" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_1\:Retrieved_Parameter_8\:description = "no parameter defined" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_1\:Retrieved_Parameter_9\:name = "not used" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_1\:Retrieved_Parameter_9\:unit = "none" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_1\:Retrieved_Parameter_9\:description = "no parameter defined" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_2\:Retrieved_Parameter_0\:name = "SSS" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_2\:Retrieved_Parameter_0\:unit = "Practical Salinity Unit (PSU)" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_2\:Retrieved_Parameter_0\:description = "Surface salinity of the sea at gridpoint" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_2\:Retrieved_Parameter_1\:name = "SST" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_2\:Retrieved_Parameter_1\:unit = "Kelvin" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_2\:Retrieved_Parameter_1\:description = "Surface temperature of the sea at gridpoint" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_2\:Retrieved_Parameter_2\:name = "UN10" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_2\:Retrieved_Parameter_2\:unit = "m.s-1" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_2\:Retrieved_Parameter_2\:description = "U component of neutral wind 10m above surface" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_2\:Retrieved_Parameter_3\:name = "VN10" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_2\:Retrieved_Parameter_3\:unit = "m.s-1" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_2\:Retrieved_Parameter_3\:description = "V component of neutral wind 10m above surface" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_2\:Retrieved_Parameter_4\:name = "tec" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_2\:Retrieved_Parameter_4\:unit = "tecu" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_2\:Retrieved_Parameter_4\:description = "Total Electronic Content of the ionosphere below SMOS" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_2\:Retrieved_Parameter_5\:name = "not used" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_2\:Retrieved_Parameter_5\:unit = "none" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_2\:Retrieved_Parameter_5\:description = "no parameter defined" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_2\:Retrieved_Parameter_6\:name = "not used" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_2\:Retrieved_Parameter_6\:unit = "none" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_2\:Retrieved_Parameter_6\:description = "no parameter defined" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_2\:Retrieved_Parameter_7\:name = "not used" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_2\:Retrieved_Parameter_7\:unit = "none" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_2\:Retrieved_Parameter_7\:description = "no parameter defined" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_2\:Retrieved_Parameter_8\:name = "not used" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_2\:Retrieved_Parameter_8\:unit = "none" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_2\:Retrieved_Parameter_8\:description = "no parameter defined" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_2\:Retrieved_Parameter_9\:name = "not used" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_2\:Retrieved_Parameter_9\:unit = "none" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_2\:Retrieved_Parameter_9\:description = "no parameter defined" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_3\:Retrieved_Parameter_0\:name = "Acard" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_3\:Retrieved_Parameter_0\:unit = "dl" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_3\:Retrieved_Parameter_0\:description = "Acard coefficient for cardioid model" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_3\:Retrieved_Parameter_1\:name = "SST" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_3\:Retrieved_Parameter_1\:unit = "Kelvin" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_3\:Retrieved_Parameter_1\:description = "Surface temperature of the sea at gridpoint" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_3\:Retrieved_Parameter_2\:name = "not used" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_3\:Retrieved_Parameter_2\:unit = "none" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_3\:Retrieved_Parameter_2\:description = "no parameter defined" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_3\:Retrieved_Parameter_3\:name = "not used" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_3\:Retrieved_Parameter_3\:unit = "none" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_3\:Retrieved_Parameter_3\:description = "no parameter defined" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_3\:Retrieved_Parameter_4\:name = "not used" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_3\:Retrieved_Parameter_4\:unit = "none" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_3\:Retrieved_Parameter_4\:description = "no parameter defined" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_3\:Retrieved_Parameter_5\:name = "not used" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_3\:Retrieved_Parameter_5\:unit = "none" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_3\:Retrieved_Parameter_5\:description = "no parameter defined" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_3\:Retrieved_Parameter_6\:name = "not used" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_3\:Retrieved_Parameter_6\:unit = "none" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_3\:Retrieved_Parameter_6\:description = "no parameter defined" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_3\:Retrieved_Parameter_7\:name = "not used" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_3\:Retrieved_Parameter_7\:unit = "none" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_3\:Retrieved_Parameter_7\:description = "no parameter defined" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_3\:Retrieved_Parameter_8\:name = "not used" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_3\:Retrieved_Parameter_8\:unit = "none" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_3\:Retrieved_Parameter_8\:description = "no parameter defined" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_3\:Retrieved_Parameter_9\:name = "not used" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_3\:Retrieved_Parameter_9\:unit = "none" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_3\:Retrieved_Parameter_9\:description = "no parameter defined" ;
		string :VH\:SPH\:MI\:SPH_Descriptor = "MIR_OSUDP2_SPH" ;
		string :VH\:SPH\:MI\:Checksum = "2323233818" ;
		string :VH\:SPH\:MI\:Header_Schema = "HDR_SM_XXXX_MIR_OSUDP2_0400.xsd" ;
		string :VH\:SPH\:MI\:Datablock_Schema = "DBL_SM_XXXX_MIR_OSUDP2_0401.binXschema.xml" ;
		string :VH\:SPH\:MI\:Header_Size = "168709" ;
		string :VH\:SPH\:MI\:Datablock_Size = "00020206504" ;
		string :VH\:SPH\:MI\:HW_Identifier = "0003" ;
		string :VH\:SPH\:MI\:TI\:Precise_Validity_Start = "UTC=2021-06-30T21:09:12.434579" ;
		string :VH\:SPH\:MI\:TI\:Precise_Validity_Stop = "UTC=2021-06-30T22:02:28.074411" ;
		string :VH\:SPH\:MI\:TI\:Abs_Orbit_Start = "+61281" ;
		string :VH\:SPH\:MI\:TI\:Start_Time_ANX_T = "1286.293116" ;
		string :VH\:SPH\:MI\:TI\:Abs_Orbit_Stop = "+61281" ;
		string :VH\:SPH\:MI\:TI\:Stop_Time_ANX_T = "4481.932948" ;
		string :VH\:SPH\:MI\:TI\:UTC_at_ANX = "UTC=2021-06-30T20:47:46.141463" ;
		string :VH\:SPH\:MI\:TI\:Long_at_ANX = "+138.381497" ;
		string :VH\:SPH\:MI\:TI\:Ascending_Flag = "D" ;
		string :VH\:SPH\:MI\:TI\:Polarisation_Flag = "F" ;
		string :VH\:SPH\:LODS\:Data_Set_0\:DS_Name = "SSS_SWATH" ;
		string :VH\:SPH\:LODS\:Data_Set_0\:DS_Type = "M" ;
		string :VH\:SPH\:LODS\:Data_Set_0\:DS_Size = "0020206504" ;
		string :VH\:SPH\:LODS\:Data_Set_0\:DS_Offset = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_0\:Num_DSR = "0000106350" ;
		string :VH\:SPH\:LODS\:Data_Set_0\:DSR_Size = "00000190" ;
		string :VH\:SPH\:LODS\:Data_Set_0\:Byte_Order = "0123" ;
		string :VH\:SPH\:LODS\:Data_Set_1\:DS_Name = "L1C_OS_FILE" ;
		string :VH\:SPH\:LODS\:Data_Set_1\:DS_Type = "R" ;
		string :VH\:SPH\:LODS\:Data_Set_1\:DS_Size = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_1\:DS_Offset = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_1\:Ref_Filename = "SM_OPER_MIR_SCSF1C_20210630T210913_20210630T220228_724_001_1" ;
		string :VH\:SPH\:LODS\:Data_Set_1\:Num_DSR = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_1\:DSR_Size = "00000000" ;
		string :VH\:SPH\:LODS\:Data_Set_1\:Byte_Order = "0000" ;
		string :VH\:SPH\:LODS\:Data_Set_2\:DS_Name = "DGG_FILE" ;
		string :VH\:SPH\:LODS\:Data_Set_2\:DS_Type = "R" ;
		string :VH\:SPH\:LODS\:Data_Set_2\:DS_Size = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_2\:DS_Offset = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_2\:Ref_Filename = "SM_OPER_AUX_DGG____20050101T000000_20500101T000000_300_003_3" ;
		string :VH\:SPH\:LODS\:Data_Set_2\:Num_DSR = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_2\:DSR_Size = "00000000" ;
		string :VH\:SPH\:LODS\:Data_Set_2\:Byte_Order = "0000" ;
		string :VH\:SPH\:LODS\:Data_Set_3\:DS_Name = "IERS_BULLETIN_B_FILE" ;
		string :VH\:SPH\:LODS\:Data_Set_3\:DS_Type = "R" ;
		string :VH\:SPH\:LODS\:Data_Set_3\:DS_Size = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_3\:DS_Offset = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_3\:Ref_Filename = "SM_OPER_AUX_BULL_B_20210402T000000_20500101T000000_120_001_3" ;
		string :VH\:SPH\:LODS\:Data_Set_3\:Num_DSR = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_3\:DSR_Size = "00000000" ;
		string :VH\:SPH\:LODS\:Data_Set_3\:Byte_Order = "0000" ;
		string :VH\:SPH\:LODS\:Data_Set_4\:DS_Name = "BESTFITPLANE_FILE" ;
		string :VH\:SPH\:LODS\:Data_Set_4\:DS_Type = "R" ;
		string :VH\:SPH\:LODS\:Data_Set_4\:DS_Size = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_4\:DS_Offset = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_4\:Ref_Filename = "SM_OPER_AUX_BFP____20050101T000000_20500101T000000_340_004_3" ;
		string :VH\:SPH\:LODS\:Data_Set_4\:Num_DSR = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_4\:DSR_Size = "00000000" ;
		string :VH\:SPH\:LODS\:Data_Set_4\:Byte_Order = "0000" ;
		string :VH\:SPH\:LODS\:Data_Set_5\:DS_Name = "MISPOINTING_FILE" ;
		string :VH\:SPH\:LODS\:Data_Set_5\:DS_Type = "R" ;
		string :VH\:SPH\:LODS\:Data_Set_5\:DS_Size = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_5\:DS_Offset = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_5\:Ref_Filename = "SM_OPER_AUX_MISP___20050101T000000_20500101T000000_300_004_3" ;
		string :VH\:SPH\:LODS\:Data_Set_5\:Num_DSR = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_5\:DSR_Size = "00000000" ;
		string :VH\:SPH\:LODS\:Data_Set_5\:Byte_Order = "0000" ;
		string :VH\:SPH\:LODS\:Data_Set_6\:DS_Name = "ECMWF_FILE" ;
		string :VH\:SPH\:LODS\:Data_Set_6\:DS_Type = "R" ;
		string :VH\:SPH\:LODS\:Data_Set_6\:DS_Size = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_6\:DS_Offset = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_6\:Ref_Filename = "SM_OPER_AUX_ECMWF__20210630T210900_20210630T221540_318_001_3" ;
		string :VH\:SPH\:LODS\:Data_Set_6\:Num_DSR = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_6\:DSR_Size = "00000000" ;
		string :VH\:SPH\:LODS\:Data_Set_6\:Byte_Order = "0000" ;
		string :VH\:SPH\:LODS\:Data_Set_7\:DS_Name = "FLAT_SEA_FILE" ;
		string :VH\:SPH\:LODS\:Data_Set_7\:DS_Type = "R" ;
		string :VH\:SPH\:LODS\:Data_Set_7\:DS_Size = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_7\:DS_Offset = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_7\:Ref_Filename = "SM_OPER_AUX_FLTSEA_20050101T000000_20500101T000000_001_012_3" ;
		string :VH\:SPH\:LODS\:Data_Set_7\:Num_DSR = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_7\:DSR_Size = "00000000" ;
		string :VH\:SPH\:LODS\:Data_Set_7\:Byte_Order = "0000" ;
		string :VH\:SPH\:LODS\:Data_Set_8\:DS_Name = "ROUGHNESS_IPSL_FILE" ;
		string :VH\:SPH\:LODS\:Data_Set_8\:DS_Type = "R" ;
		string :VH\:SPH\:LODS\:Data_Set_8\:DS_Size = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_8\:DS_Offset = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_8\:Ref_Filename = "SM_OPER_AUX_RGHNS1_20050101T000000_20500101T000000_001_016_3" ;
		string :VH\:SPH\:LODS\:Data_Set_8\:Num_DSR = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_8\:DSR_Size = "00000000" ;
		string :VH\:SPH\:LODS\:Data_Set_8\:Byte_Order = "0000" ;
		string :VH\:SPH\:LODS\:Data_Set_9\:DS_Name = "ROUGHNESS_IFREMER_FILE" ;
		string :VH\:SPH\:LODS\:Data_Set_9\:DS_Type = "R" ;
		string :VH\:SPH\:LODS\:Data_Set_9\:DS_Size = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_9\:DS_Offset = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_9\:Ref_Filename = "SM_OPER_AUX_RGHNS2_20050101T000000_20500101T000000_001_013_3" ;
		string :VH\:SPH\:LODS\:Data_Set_9\:Num_DSR = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_9\:DSR_Size = "00000000" ;
		string :VH\:SPH\:LODS\:Data_Set_9\:Byte_Order = "0000" ;
		string :VH\:SPH\:LODS\:Data_Set_10\:DS_Name = "ROUGHNESS_ICM_CSIC_FILE" ;
		string :VH\:SPH\:LODS\:Data_Set_10\:DS_Type = "R" ;
		string :VH\:SPH\:LODS\:Data_Set_10\:DS_Size = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_10\:DS_Offset = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_10\:Ref_Filename = "SM_OPER_AUX_RGHNS3_20050101T000000_20500101T000000_001_016_3" ;
		string :VH\:SPH\:LODS\:Data_Set_10\:Num_DSR = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_10\:DSR_Size = "00000000" ;
		string :VH\:SPH\:LODS\:Data_Set_10\:Byte_Order = "0000" ;
		string :VH\:SPH\:LODS\:Data_Set_11\:DS_Name = "GALAXY_OS_FILE" ;
		string :VH\:SPH\:LODS\:Data_Set_11\:DS_Type = "R" ;
		string :VH\:SPH\:LODS\:Data_Set_11\:DS_Size = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_11\:DS_Offset = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_11\:Ref_Filename = "SM_OPER_AUX_GAL_OS_20050101T000000_20500101T000000_001_011_3" ;
		string :VH\:SPH\:LODS\:Data_Set_11\:Num_DSR = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_11\:DSR_Size = "00000000" ;
		string :VH\:SPH\:LODS\:Data_Set_11\:Byte_Order = "0000" ;
		string :VH\:SPH\:LODS\:Data_Set_12\:DS_Name = "GALAXY_2OS_FILE" ;
		string :VH\:SPH\:LODS\:Data_Set_12\:DS_Type = "R" ;
		string :VH\:SPH\:LODS\:Data_Set_12\:DS_Size = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_12\:DS_Offset = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_12\:Ref_Filename = "SM_OPER_AUX_GAL2OS_20050101T000000_20500101T000000_001_016_3" ;
		string :VH\:SPH\:LODS\:Data_Set_12\:Num_DSR = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_12\:DSR_Size = "00000000" ;
		string :VH\:SPH\:LODS\:Data_Set_12\:Byte_Order = "0000" ;
		string :VH\:SPH\:LODS\:Data_Set_13\:DS_Name = "SUNGLINT_FILE" ;
		string :VH\:SPH\:LODS\:Data_Set_13\:DS_Type = "R" ;
		string :VH\:SPH\:LODS\:Data_Set_13\:DS_Size = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_13\:DS_Offset = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_13\:Ref_Filename = "SM_OPER_AUX_SGLINT_20050101T000000_20500101T000000_001_012_3" ;
		string :VH\:SPH\:LODS\:Data_Set_13\:Num_DSR = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_13\:DSR_Size = "00000000" ;
		string :VH\:SPH\:LODS\:Data_Set_13\:Byte_Order = "0000" ;
		string :VH\:SPH\:LODS\:Data_Set_14\:DS_Name = "ATMOS_FILE" ;
		string :VH\:SPH\:LODS\:Data_Set_14\:DS_Type = "R" ;
		string :VH\:SPH\:LODS\:Data_Set_14\:DS_Size = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_14\:DS_Offset = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_14\:Ref_Filename = "SM_OPER_AUX_ATMOS__20050101T000000_20500101T000000_001_010_3" ;
		string :VH\:SPH\:LODS\:Data_Set_14\:Num_DSR = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_14\:DSR_Size = "00000000" ;
		string :VH\:SPH\:LODS\:Data_Set_14\:Byte_Order = "0000" ;
		string :VH\:SPH\:LODS\:Data_Set_15\:DS_Name = "DISTAN_FILE" ;
		string :VH\:SPH\:LODS\:Data_Set_15\:DS_Type = "R" ;
		string :VH\:SPH\:LODS\:Data_Set_15\:DS_Size = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_15\:DS_Offset = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_15\:Ref_Filename = "SM_OPER_AUX_DISTAN_20050101T000000_20500101T000000_001_011_3" ;
		string :VH\:SPH\:LODS\:Data_Set_15\:Num_DSR = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_15\:DSR_Size = "00000000" ;
		string :VH\:SPH\:LODS\:Data_Set_15\:Byte_Order = "0000" ;
		string :VH\:SPH\:LODS\:Data_Set_16\:DS_Name = "CLIMATOLOGY_SSS_FILE" ;
		string :VH\:SPH\:LODS\:Data_Set_16\:DS_Type = "R" ;
		string :VH\:SPH\:LODS\:Data_Set_16\:DS_Size = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_16\:DS_Offset = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_16\:Ref_Filename = "SM_OPER_AUX_SSS____20050101T000000_20500101T000000_001_014_3" ;
		string :VH\:SPH\:LODS\:Data_Set_16\:Num_DSR = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_16\:DSR_Size = "00000000" ;
		string :VH\:SPH\:LODS\:Data_Set_16\:Byte_Order = "0000" ;
		string :VH\:SPH\:LODS\:Data_Set_17\:DS_Name = "CLIMATOLOGY_SSSCLI_FILE" ;
		string :VH\:SPH\:LODS\:Data_Set_17\:DS_Type = "R" ;
		string :VH\:SPH\:LODS\:Data_Set_17\:DS_Size = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_17\:DS_Offset = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_17\:Ref_Filename = "SM_OPER_AUX_SSSCLI_20050101T000000_20500101T000000_001_002_3" ;
		string :VH\:SPH\:LODS\:Data_Set_17\:Num_DSR = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_17\:DSR_Size = "00000000" ;
		string :VH\:SPH\:LODS\:Data_Set_17\:Byte_Order = "0000" ;
		string :VH\:SPH\:LODS\:Data_Set_18\:DS_Name = "OCEAN_SALINITY_CONFIG_FILE" ;
		string :VH\:SPH\:LODS\:Data_Set_18\:DS_Type = "R" ;
		string :VH\:SPH\:LODS\:Data_Set_18\:DS_Size = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_18\:DS_Offset = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_18\:Ref_Filename = "SM_OPER_AUX_CNFOSF_20050101T000000_20500101T000000_001_032_3" ;
		string :VH\:SPH\:LODS\:Data_Set_18\:Num_DSR = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_18\:DSR_Size = "00000000" ;
		string :VH\:SPH\:LODS\:Data_Set_18\:Byte_Order = "0000" ;
		string :VH\:SPH\:LODS\:Data_Set_19\:DS_Name = "OTT1F_FILE" ;
		string :VH\:SPH\:LODS\:Data_Set_19\:DS_Type = "R" ;
		string :VH\:SPH\:LODS\:Data_Set_19\:DS_Size = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_19\:DS_Offset = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_19\:Ref_Filename = "SM_OPER_AUX_OTT1F__20210624T082406_20500101T000000_700_001_1" ;
		string :VH\:SPH\:LODS\:Data_Set_19\:Num_DSR = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_19\:DSR_Size = "00000000" ;
		string :VH\:SPH\:LODS\:Data_Set_19\:Byte_Order = "0000" ;
		string :VH\:SPH\:LODS\:Data_Set_20\:DS_Name = "OTT2F_FILE" ;
		string :VH\:SPH\:LODS\:Data_Set_20\:DS_Type = "R" ;
		string :VH\:SPH\:LODS\:Data_Set_20\:DS_Size = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_20\:DS_Offset = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_20\:Ref_Filename = "SM_OPER_AUX_OTT2F__20210624T082406_20500101T000000_700_001_1" ;
		string :VH\:SPH\:LODS\:Data_Set_20\:Num_DSR = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_20\:DSR_Size = "00000000" ;
		string :VH\:SPH\:LODS\:Data_Set_20\:Byte_Order = "0000" ;
		string :VH\:SPH\:LODS\:Data_Set_21\:DS_Name = "OTT3F_FILE" ;
		string :VH\:SPH\:LODS\:Data_Set_21\:DS_Type = "R" ;
		string :VH\:SPH\:LODS\:Data_Set_21\:DS_Size = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_21\:DS_Offset = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_21\:Ref_Filename = "SM_OPER_AUX_OTT3F__20210624T082406_20500101T000000_700_001_1" ;
		string :VH\:SPH\:LODS\:Data_Set_21\:Num_DSR = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_21\:DSR_Size = "00000000" ;
		string :VH\:SPH\:LODS\:Data_Set_21\:Byte_Order = "0000" ;
		string :VH\:SPH\:LODS\:Data_Set_22\:DS_Name = "DGGRFI_FILE" ;
		string :VH\:SPH\:LODS\:Data_Set_22\:DS_Type = "R" ;
		string :VH\:SPH\:LODS\:Data_Set_22\:DS_Size = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_22\:DS_Offset = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_22\:Ref_Filename = "SM_OPER_AUX_DGGRFI_20210629T000711_20500101T000000_600_001_1" ;
		string :VH\:SPH\:LODS\:Data_Set_22\:Num_DSR = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_22\:DSR_Size = "00000000" ;
		string :VH\:SPH\:LODS\:Data_Set_22\:Byte_Order = "0000" ;
		string :VH\:SPH\:LODS\:Data_Set_23\:DS_Name = "MIXED_SCENE_OTT_FILE" ;
		string :VH\:SPH\:LODS\:Data_Set_23\:DS_Type = "R" ;
		string :VH\:SPH\:LODS\:Data_Set_23\:DS_Size = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_23\:DS_Offset = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_23\:Ref_Filename = "SM_OPER_AUX_MSOTT__20050101T000000_20500101T000000_001_002_3" ;
		string :VH\:SPH\:LODS\:Data_Set_23\:Num_DSR = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_23\:DSR_Size = "00000000" ;
		string :VH\:SPH\:LODS\:Data_Set_23\:Byte_Order = "0000" ;
		string :VH\:SPH\:L2PL\:Start_Lat = "+075.719335" ;
		string :VH\:SPH\:L2PL\:Start_Long = "+097.548779" ;
		string :VH\:SPH\:L2PL\:Stop_Lat = "-081.598965" ;
		string :VH\:SPH\:L2PL\:Stop_Long = "-150.028234" ;
		string :VH\:SPH\:L2PL\:Mid_Lat = "+005.419643" ;
		string :VH\:SPH\:L2PL\:Mid_Lon = "-052.859901" ;
		string :VH\:SPH\:L2PL\:Southernmost_Latitude = "-067.069000" ;
		string :VH\:SPH\:L2PL\:Southernmost_Gridpoint_ID = "6166549" ;
		string :VH\:SPH\:L2PL\:Northernmost_Latitude = "+079.646004" ;
		string :VH\:SPH\:L2PL\:Northernmost_Gridpoint_ID = "0002902" ;
		string :VH\:SPH\:L2PL\:Easternmost_Longitude = "+049.222000" ;
		string :VH\:SPH\:L2PL\:Easternmost_Gridpoint_ID = "4084941" ;
		string :VH\:SPH\:L2PL\:Westernmost_Longitude = "-090.652000" ;
		string :VH\:SPH\:L2PL\:Westernmost_Gridpoint_ID = "6155252" ;
		string :VH\:MPH\:Ref_Doc = "SO-TN-IDR-GS-0006" ;
		string :VH\:MPH\:Acquisition_Station = "SVLD" ;
		string :VH\:MPH\:Processing_Centre = "ESAC" ;
		string :VH\:MPH\:Logical_Proc_Centre = "FPC" ;
		string :VH\:MPH\:Product_Confidence = "NOMINAL" ;
		string :VH\:MPH\:OI\:Phase = "+001" ;
		string :VH\:MPH\:OI\:Cycle = "+037" ;
		string :VH\:MPH\:OI\:Rel_Orbit = "+01161" ;
		string :VH\:MPH\:OI\:Abs_Orbit = "+61281" ;
		string :VH\:MPH\:OI\:OSV_TAI = "TAI=2021-06-30T21:08:37.000000" ;
		string :VH\:MPH\:OI\:OSV_UTC = "UTC=2021-06-30T21:08:00.000000" ;
		string :VH\:MPH\:OI\:OSV_UT1 = "UT1=2021-06-30T21:08:00.590000" ;
		string :VH\:MPH\:OI\:X_Position = "-0616039.695" ;
		string :VH\:MPH\:OI\:Y_Position = "+2121521.304" ;
		string :VH\:MPH\:OI\:Z_Position = "+6778739.127" ;
		string :VH\:MPH\:OI\:X_Velocity = "+5304.621980" ;
		string :VH\:MPH\:OI\:Y_Velocity = "-4977.113140" ;
		string :VH\:MPH\:OI\:Z_Velocity = "+2035.575410" ;
		string :VH\:MPH\:OI\:Vector_Source = "FP" ;
		:history = "Mon Oct  2 16:01:51 2023: ncks -d n_grid_points,100,92700,1800 -v SSS_corr,Sigma_SSS_corr,Latitude,Longitude,Mean_acq_time,Dg_quality_SSS_corr /scratch1/NCEPDEV/stmp4/Shastri.Paturi/forAndrew/gdas.20210701/00/SSS/SM_OPER_MIR_OSUDP2_20210630T210913_20210630T220228_700_001_1.nc sss_smos_1_sub.nc" ;
		:NCO = "netCDF Operators version 5.0.6 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco)" ;
data:

 Dg_quality_SSS_corr = _, _, _, _, _, _, _, _, _, 426, _, _, _, _, _, _, 70, 
    76, 157, 226, 369, _, 397, 77, 56, 105, 162, _, 78, 57, _, _, 185, _, _, 
    161, 164, _, _, _, _, _, _, _, _, _, _, _, _, _, 186, 447 ;

 Latitude = 84.474, 79.093, 79.069, 85.988, 73.646, 74.369, 73.373, 68.824, 
    67.431, 67.911, 61.056, 66.861, 64.861, 63.581, 61.064, 49.872, 48.513, 
    46.599, 43.993, 46.536, 47.555, 46.194, 43.333, 32.862, 31.318, 28.788, 
    32.755, 32.526, 21.871, 20.343, 17.874, 15.329, 20.809, 10.47, 9.402, 
    11.548, 11.246, 0.365, -1.881, -31.722, -34.284, -36.43, -45.173, 
    -49.272, -49.917, -52.05, -54.981, -47.587, -52.566, -60.212, -62.353, 
    -64.333 ;

 Longitude = 9.96, -6.847, 15.206, 21.943, -7.968, -26.325, 8.154, -21.809, 
    -35.023, -11.93, -30.459, -41.569, -43.384, -46.592, -46.251, -37.368, 
    -40.068, -42.775, -46.637, -35.473, -49.166, -51.088, -50.423, -44.497, 
    -47.041, -50.208, -50.903, -53, -47.445, -49.855, -52.654, -53.977, 
    -54.428, -49.443, -52.964, -47.409, -55.798, -50.84, -52.914, -58.202, 
    -56.971, -55.46, -69.335, -63.251, -71.935, -68.916, -67.195, -75.662, 
    -58.381, -78.897, -76.082, -86.052 ;

 Mean_acq_time = 7851.884, 7851.884, _, 7851.883, 7851.885, _, 7851.885, 
    7851.886, _, 7851.887, 7851.888, _, _, _, 7851.889, 7851.89, 7851.891, 
    7851.891, 7851.892, 7851.891, 7851.892, 7851.892, 7851.893, 7851.894, 
    7851.894, 7851.895, 7851.895, 7851.895, 7851.896, 7851.896, 7851.896, 
    7851.897, 7851.896, 7851.898, 7851.898, 7851.898, 7851.898, _, _, _, _, 
    7851.907, _, 7851.91, _, _, _, 7851.91, 7851.911, 7851.912, 7851.913, 
    7851.914 ;

 SSS_corr = _, _, _, _, 28.72996, _, _, 32.20172, _, 34.32167, 33.84064, _, 
    _, _, _, 34.39512, 34.14527, 33.85896, 32.81892, 37.6133, 33.1171, _, 
    31.79991, 36.53445, 38.26277, 37.38822, 36.66851, _, 38.08805, 37.35236, 
    35.68861, 32.68691, 35.8759, 36.5416, 31.50342, 34.18812, 32.44438, _, _, 
    _, _, _, _, 34.83915, _, _, _, _, _, 33.43178, 34.17802, 31.58817 ;

 Sigma_SSS_corr = _, _, _, _, 2.255848, _, _, 3.373118, _, 4.289972, 
    0.966469, _, _, _, _, 0.7200613, 0.9667612, 1.166589, 0.862876, 1.606015, 
    3.603568, _, 3.201073, 0.5792597, 0.508775, 0.6778937, 1.006906, _, 
    0.7903381, 0.6655976, 0.7761204, 1.059877, 1.433936, 0.7581352, 
    0.5698198, 1.306699, 1.07838, _, _, _, _, _, _, 1.56893, _, _, _, _, _, 
    2.569222, 2.849992, 3.374218 ;
}
