netcdf output_2 {
dimensions:
	Rows = 15 ;
	Columns = 50 ;
variables:
	float IceConc(Rows, Columns) ;
		IceConc:_FillValue = -999.f ;
		IceConc:coordinates = "Longitude Latitude" ;
		IceConc:long_name = "Ice Concentration" ;
		IceConc:units = "%" ;
		IceConc:valid_range = 0.f, 100.f ;
	byte IceMap(Rows, Columns) ;
		IceMap:_FillValue = -3b ;
		IceMap:coordinates = "Longitude Latitude" ;
		IceMap:long_name = "Ice Cover map codes" ;
		IceMap:units = "1" ;
		IceMap:valid_range = -2b, 2b ;
	float IceRetrPct ;
		IceRetrPct:long_name = "% of valid ice cover and concentration retrievals of all water pixels" ;
		IceRetrPct:units = "%" ;
		IceRetrPct:_FillValue = 0.f ;
		IceRetrPct:valid_range = 0.f, 100.f ;
	float IceSrfTemp(Rows, Columns) ;
		IceSrfTemp:_FillValue = -999.f ;
		IceSrfTemp:coordinates = "Longitude Latitude" ;
		IceSrfTemp:long_name = "Ice Surface Temp" ;
		IceSrfTemp:units = "Kelvin(K)" ;
		IceSrfTemp:valid_range = 100.f, 390.f ;
	float IceTermntPct ;
		IceTermntPct:long_name = "% of terminated ice cover and concentration retrievals of all processed pixels" ;
		IceTermntPct:units = "%" ;
		IceTermntPct:_FillValue = 0.f ;
		IceTermntPct:valid_range = 0.f, 100.f ;
	float Latitude(Rows, Columns) ;
		Latitude:long_name = "Latitude" ;
		Latitude:_FillValue = -999.f ;
		Latitude:units = "degrees_north" ;
		Latitude:valid_range = -90.f, 90.f ;
		Latitude:comments = "Pixel latitude in field Latitude (degree)" ;
	float Longitude(Rows, Columns) ;
		Longitude:long_name = "Longitude" ;
		Longitude:_FillValue = -999.f ;
		Longitude:units = "degrees_east" ;
		Longitude:valid_range = -180.f, 180.f ;
		Longitude:comments = "Pixel longitude in field Longitude (degree)" ;
	float MaxIceConc ;
		MaxIceConc:long_name = "Max ice concentration retrieval" ;
		MaxIceConc:_FillValue = -999.f ;
		MaxIceConc:units = "%" ;
	float MeanIceConc ;
		MeanIceConc:long_name = "Mean ice concentration retrieval" ;
		MeanIceConc:_FillValue = -999.f ;
		MeanIceConc:units = "%" ;
	float MinIceConc ;
		MinIceConc:long_name = "Min ice concentration retrieval" ;
		MinIceConc:_FillValue = -999.f ;
		MinIceConc:units = "%" ;
	byte NumOfQACategories ;
		NumOfQACategories:long_name = "Number of QA flag values" ;
		NumOfQACategories:_FillValue = -128b ;
		NumOfQACategories:units = "1" ;
	int QCFlags(Rows, Columns) ;
		QCFlags:_FillValue = -1 ;
		QCFlags:coordinates = "Longitude Latitude" ;
		QCFlags:long_name = "QCFlags" ;
		QCFlags:units = "1" ;
	float STDIceConc ;
		STDIceConc:long_name = "Standard deviation of ice concentration retrievals" ;
		STDIceConc:_FillValue = -999.f ;
		STDIceConc:units = "%" ;
	byte SearchWindowSize ;
		SearchWindowSize:long_name = "Pixel size of search window to determine tie-point" ;
		SearchWindowSize:_FillValue = -128b ;
		SearchWindowSize:units = "1" ;
	int StartColumn ;
		StartColumn:long_name = "Start column index" ;
		StartColumn:units = "1" ;
	int StartRow ;
		StartRow:long_name = "Start row index" ;
		StartRow:units = "1" ;
	byte SummaryQC_Ice_Concentration(Rows, Columns) ;
		SummaryQC_Ice_Concentration:_FillValue = -128b ;
		SummaryQC_Ice_Concentration:coordinates = "Longitude Latitude" ;
		SummaryQC_Ice_Concentration:long_name = "User-level summary QC: 0=Normal, 1=Uncertain, 2=Non-Retrievable, 3=Bad" ;
		SummaryQC_Ice_Concentration:units = "1" ;
		SummaryQC_Ice_Concentration:valid_range = 0b, 3b ;
	int TotDaytimePixs ;
		TotDaytimePixs:long_name = "Total number of daytime valid retrievals" ;
		TotDaytimePixs:_FillValue = 0 ;
		TotDaytimePixs:units = "1" ;
	int TotIceRetrvls ;
		TotIceRetrvls:long_name = "Total number of valid ice cover and concentration retrievals" ;
		TotIceRetrvls:_FillValue = 0 ;
		TotIceRetrvls:units = "1" ;
	int TotIceTermnt ;
		TotIceTermnt:long_name = "Total number of terminated ice cover and concentration retrievals" ;
		TotIceTermnt:_FillValue = 0 ;
		TotIceTermnt:units = "1" ;
	int TotNighttimePixs ;
		TotNighttimePixs:long_name = "Total number of nighttime valid retrievals" ;
		TotNighttimePixs:_FillValue = 0 ;
		TotNighttimePixs:units = "1" ;
	int TotWaterPixs ;
		TotWaterPixs:long_name = "Total number of pixels w. water surface" ;
		TotWaterPixs:_FillValue = 0 ;
		TotWaterPixs:units = "1" ;
	int Tot_QA_BadData ;
		Tot_QA_BadData:long_name = "Total number of pixels with QA category 4 (Bad data)" ;
		Tot_QA_BadData:_FillValue = 0 ;
		Tot_QA_BadData:units = "1" ;
	int Tot_QA_Nonretrievable ;
		Tot_QA_Nonretrievable:long_name = "Total number of pixels with QA category 3 (Non-retrievable)" ;
		Tot_QA_Nonretrievable:_FillValue = 0 ;
		Tot_QA_Nonretrievable:units = "1" ;
	int Tot_QA_Normal ;
		Tot_QA_Normal:long_name = "Total number of pixels with QA category 1 (Normal of optimal)" ;
		Tot_QA_Normal:_FillValue = 0 ;
		Tot_QA_Normal:units = "1" ;
	int Tot_QA_Uncertain ;
		Tot_QA_Uncertain:long_name = "Total number of pixels with QA category 2 (Uncertain or suboptimal)" ;
		Tot_QA_Uncertain:_FillValue = 0 ;
		Tot_QA_Uncertain:units = "1" ;

// global attributes:
		:Conventions = "CF-1.6,ACDD 1.3" ;
		:Metadata_Conventions = "CF-1.6, Unidata Dataset Discovery v1.0" ;
		:standard_name_vocabulary = "CF Standard Name Table v76" ;
		:institution = "DOC/NOAA/NESDIS/OSPO > Office of Satellite and Product Operations, NESDIS, NOAA, U.S. Department of Commerce." ;
		:naming_authority = "gov.noaa.nesdis.ncei." ;
		:processing_level = "NOAA Level 2" ;
		:production_site = "NCCF" ;
		:production_environment = "prod" ;
		:sensor_band_identifier = "M3,M5,M7,M10,M15,M16" ;
		:sensor_band_central_radiation_wavelength = "0.488um,0.672um,0.865um,1.61um,10.763um,12.013um" ;
		:satellite_name = "NOAA-20" ;
		:instrument = "VIIRS" ;
		:project = "NESDIS Common Cloud Framework" ;
		:summary = "Enterprise Ice Concentration/ Ice Mask/ Ice Surface Temperature Products" ;
		:history = "Tue Aug 20 14:35:27 2024: ncks -d Columns,902,1000,2 -d Rows,422,451,2 JRR-IceConcentration_v3r3_j01_s202406180952557_e202406180954184_c202406181023196.nc output_2.nc\nEnterprise Ice Concentration Algorithm v1.1.0" ;
		:references = "N/A" ;
		:resolution = "750M" ;
		:time_coverage_start = "2024-06-18T09:52:55Z" ;
		:time_coverage_end = "2024-06-18T09:54:18Z" ;
		:date_created = "2024-06-18T10:23:19Z" ;
		:geospatial_lat_units = "degrees_north" ;
		:geospatial_lon_units = "degrees_east" ;
		:publisher_name = "DOC/NOAA/NESDIS/OSPO > Office of Satellite and Product Operations, NESDIS, NOAA, U.S. Department of Commerce." ;
		:publisher_email = "espcoperations@noaa.gov" ;
		:publisher_url = "http://www.ospo.noaa.gov" ;
		:creator_email = "jkey@ssec.wisc.edu" ;
		:creator_name = "DOC/NOAA/NESDIS/STAR > Cryosphere Team, Center for Satellite Applications and Research, NESDIS, NOAA, U.S. Department of Commerce" ;
		:creator_url = "http://www.star.nesdis.noaa.gov" ;
		:source = "L1b data, JRR-CloudMask, JRR-CloudHeight" ;
		:keywords = "EARTH SCIENCE, CRYOSPHERE, SEA ICE, SEA ICE CONCENTRATION, ICE FRACTION, ICE EXTENT, ICE EDGES" ;
		:cdm_data_type = "Swath" ;
		:platform = "NOAA-20" ;
		:title = "JRR_IceConcentration" ;
		:metadata_link = "JRR-IceConcentration_v3r3_j01_s202406180952557_e202406180954184_c202406181023196.nc" ;
		:history_package = "Delivery Package v3r3" ;
		:product_version = "v3r3" ;
		:keywords_vocabulary = "NASA Global Change Master Directory (GCMD) Science Keywords" ;
		:geospatial_lat_max = 90.f ;
		:geospatial_lat_min = -90.f ;
		:geospatial_lat_resolution = "750 meters" ;
		:geospatial_lon_max = 180.f ;
		:geospatial_lon_min = -180.f ;
		:geospatial_lon_resolution = "750 meters" ;
		:id = "b8b29146-2936-461e-b20a-b9cf98790cbf" ;
		:geospatial_bounds = "POLYGON((66.674118 64.1376266, 12.215044 56.018959, 5.55829859 59.631855, 68.5783844 68.9835892, 66.674118 64.1376266))" ;
		:day_night_data_flag = "day" ;
		:start_orbit_number = 34108 ;
		:end_orbit_number = 34108 ;
		:ascend_descend_data_flag = 0 ;
		:geospatial_first_scanline_first_fov_lat = 64.13763f ;
		:geospatial_first_scanline_last_fov_lat = 68.98359f ;
		:geospatial_last_scanline_first_fov_lat = 56.01896f ;
		:geospatial_last_scanline_last_fov_lat = 59.63186f ;
		:geospatial_first_scanline_first_fov_lon = 66.67412f ;
		:geospatial_first_scanline_last_fov_lon = 68.57838f ;
		:geospatial_last_scanline_first_fov_lon = 12.21504f ;
		:geospatial_last_scanline_last_fov_lon = 5.558299f ;
		:NCO = "netCDF Operators version 5.0.6 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco)" ;
data:

 IceConc =
  98.34166, 92.57914, 100, 100, _, 92.13963, 100, 100, 100, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _,
  100, 100, 100, _, 100, 100, 100, 100, 100, 100, 100, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  _, _, _, 100, 100, _, 100, 100, 100, 100, 100, 100, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  _, _, _, _, 100, _, _, _, _, 100, 100, _, 100, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  _, _, _, _, 100, 89.48627, _, 98.89512, _, 100, 100, 100, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  _, _, _, 100, 100, 84.68418, _, 77.50546, _, 100, 100, 100, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _,
  100, _, _, _, 100, 86.11667, 93.27911, 100, _, 100, 100, 100, 100, _, 100, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _,
  _, 71.43365, 96.33943, _, _, 83.95166, _, 100, _, 100, _, 100, 100, 100, 
    100, 100, 98.03237, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  94.22326, 100, 100, 85.10742, _, _, 100, 100, 100, 86.36085, _, _, 100, 
    100, 100, 100, 100, 76.49621, 44.59078, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  85.69344, 91.635, 88.16773, 100, 100, _, 100, 100, _, _, _, _, _, 100, 
    99.10674, 100, 100, 100, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  100, 100, 100, 100, 100, 75.4544, 100, _, 100, 83.1703, _, _, 57.75991, 
    93.47446, 100, 72.29642, _, 83.43076, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  92.31869, 89.60022, 100, 100, 100, 100, 100, _, _, 100, _, 47.09764, _, _, 
    48.18828, 55.38328, 69.85468, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  100, 100, 100, 97.60914, 95.65573, _, _, 71.58017, 70.78253, 100, 40.73283, 
    52.17646, 53.28339, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  100, 100, 100, 100, 90.26763, _, 74.51026, 81.88432, 96.97428, 96.958, 
    43.06062, 52.76248, 43.79315, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  100, 100, 100, 99.22068, 100, 100, 72.88243, 72.11736, 57.14133, 74.96605, 
    48.98592, _, 42.24671, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 IceMap =
  1, 1, 1, 1, -2, 1, 1, 1, 1, _, _, 0, -2, _, 0, 0, 0, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -2, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1,
  1, 1, 1, -2, 1, 1, 1, 1, 1, 1, 1, _, 0, -2, _, 0, -2, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1,
  -2, 0, -2, 1, 1, 0, 1, 1, 1, 1, 1, 1, -2, -2, _, 0, -2, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1,
  0, 0, 0, 0, 1, _, -2, -2, -2, 1, 1, _, 1, -2, -2, 0, 0, 0, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1,
  0, -2, -2, 0, 1, 1, -2, 1, -2, 1, 1, 1, _, -2, -2, -2, _, _, -2, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1,
  0, 0, 0, 1, 1, 1, -2, 1, -2, 1, 1, 1, _, -2, -2, -2, 0, 0, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1,
  1, 0, 0, 0, 1, 1, 1, 1, -2, 1, 1, 1, 1, -2, 1, -2, 0, 0, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1,
  _, 1, 1, _, 0, 1, -2, 1, -2, 1, -2, 1, 1, 1, 1, 1, 1, -2, _, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1,
  1, 1, 1, 1, _, 0, 1, 1, 1, 1, -2, -2, 1, 1, 1, 1, 1, 1, 1, 0, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1,
  1, 1, 1, 1, 1, _, 1, 1, 0, 0, -2, -2, -2, 1, 1, 1, 1, 1, -2, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -2, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1,
  1, 1, 1, 1, 1, 1, 1, _, 1, 1, -2, 0, 1, 1, 1, 1, -2, 1, -2, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1,
  1, 1, 1, 1, 1, 1, 1, _, _, 1, _, 1, -2, -2, 1, 1, 1, -2, 0, 0, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1,
  1, 1, 1, 1, 1, 0, _, 1, 1, 1, 1, 1, 1, 0, 0, -2, _, -2, -2, -2, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -2, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1,
  1, 1, 1, 1, 1, 0, 1, 1, 1, 1, 1, 1, 1, -2, 0, -2, _, -2, -2, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, -2, 1, 0, 0, 0, _, -2, -2, -2, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -2, -2, 
    -1, -2, -1, -1, -1, -1, -1, -1, -1 ;

 IceRetrPct = 5.886314 ;

 IceSrfTemp =
  274.9209, 274.8062, 274.9214, 274.7943, _, 274.665, 274.5973, 274.4221, 
    274.4603, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  274.8839, 274.9639, 274.973, _, 274.7099, 274.8377, 274.6533, 274.5237, 
    274.4453, 274.4314, 274.6646, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, 274.7484, 274.8216, _, 274.8814, 274.5321, 274.5942, 274.8002, 
    274.8478, 274.6158, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, 274.6919, _, _, _, _, 274.9737, 274.7827, _, 274.6674, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, 274.8948, 274.651, _, 274.8407, _, 274.6422, 274.7932, 
    274.6945, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, 274.7605, 274.6727, 274.6691, _, 274.7073, _, 274.5918, 274.5064, 
    274.3907, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  274.7585, _, _, _, 274.6302, 274.7849, 274.9124, 274.6997, _, 274.7486, 
    274.7006, 274.4442, 274.6088, _, 274.6678, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 274.9928, 274.8151, _, _, 274.9085, _, 274.8958, _, 274.8481, _, 
    274.5542, 274.5204, 274.8527, 274.6447, 274.6751, 274.5598, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  274.3351, 274.1571, 273.9791, 273.6346, _, _, 274.7652, 274.8819, 274.5946, 
    274.8276, _, _, 274.6264, 274.7227, 274.9106, 274.631, 274.7617, 
    274.9178, 274.7668, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  273.7129, 273.8175, 274.0147, 273.0873, 273.9924, _, 274.8008, 274.757, _, 
    _, _, _, _, 274.5397, 274.9979, 274.8029, 274.8488, 274.6307, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  273.3674, 273.1697, 273.3668, 272.9165, 273.2345, 273.8546, 274.9253, _, 
    274.7198, 274.7643, _, _, 274.6973, 274.9601, 273.6242, 274.2138, _, 
    274.8115, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _,
  273.7788, 273.5576, 273.6622, 273.6536, 273.5914, 273.2065, 273.1289, _, _, 
    274.2018, _, 274.1711, _, _, 274.4727, 273.6517, 273.9172, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  273.8614, 273.7878, 273.7272, 274.054, 274.0677, _, _, 274.4107, 274.4062, 
    273.796, 274.48, 273.7475, 274.541, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  273.7503, 273.7122, 273.7489, 273.8601, 274.3159, _, 273.7474, 274.2003, 
    274.0799, 273.5551, 274.2413, 273.4915, 274.3263, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  274.0728, 274.0887, 273.7952, 274.0573, 273.9589, 273.7769, 274.1772, 
    274.5915, 274.6418, 274.3053, 274.2776, _, 274.5207, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _ ;

 IceTermntPct = 99.72612 ;

 Latitude =
  66.94942, 66.94698, 66.94451, 66.94205, 66.93958, 66.93712, 66.93463, 
    66.93217, 66.9297, 66.9272, 66.92471, 66.92223, 66.91973, 66.91723, 
    66.91472, 66.91222, 66.90971, 66.9072, 66.90468, 66.90215, 66.89961, 
    66.89709, 66.89456, 66.89201, 66.88949, 66.88696, 66.8844, 66.88187, 
    66.87932, 66.87677, 66.8742, 66.87164, 66.86909, 66.86653, 66.86395, 
    66.8614, 66.85883, 66.85624, 66.85367, 66.85108, 66.8485, 66.84592, 
    66.84332, 66.84074, 66.83816, 66.83556, 66.83297, 66.83036, 66.82776, 
    66.82515,
  66.96622, 66.96376, 66.96128, 66.9588, 66.95631, 66.95382, 66.95133, 
    66.94884, 66.94633, 66.94383, 66.94132, 66.93882, 66.93629, 66.93378, 
    66.93126, 66.92873, 66.92621, 66.92368, 66.92115, 66.9186, 66.91606, 
    66.9135, 66.91095, 66.90839, 66.90585, 66.9033, 66.90073, 66.89816, 
    66.89559, 66.89303, 66.89045, 66.88787, 66.88531, 66.88272, 66.88013, 
    66.87756, 66.87496, 66.87238, 66.86978, 66.86718, 66.86458, 66.86198, 
    66.85937, 66.85677, 66.85416, 66.85156, 66.84894, 66.84632, 66.8437, 
    66.84108,
  66.98304, 66.98055, 66.97805, 66.97555, 66.97305, 66.97054, 66.96802, 
    66.9655, 66.96297, 66.96046, 66.95794, 66.9554, 66.95287, 66.95033, 
    66.94779, 66.94524, 66.9427, 66.94015, 66.9376, 66.93504, 66.93247, 
    66.9299, 66.92734, 66.92477, 66.92221, 66.91962, 66.91705, 66.91445, 
    66.91187, 66.9093, 66.90671, 66.90411, 66.90152, 66.89892, 66.89632, 
    66.8937, 66.89111, 66.88851, 66.88589, 66.88328, 66.88065, 66.87804, 
    66.87541, 66.8728, 66.87016, 66.86755, 66.86491, 66.86229, 66.85965, 
    66.85701,
  66.99986, 66.99734, 66.99483, 66.99229, 66.98977, 66.98724, 66.9847, 
    66.98218, 66.97964, 66.9771, 66.97455, 66.97199, 66.96944, 66.9669, 
    66.96433, 66.96176, 66.95921, 66.95663, 66.95407, 66.95148, 66.94889, 
    66.94631, 66.94373, 66.94114, 66.93855, 66.93595, 66.93336, 66.93076, 
    66.92816, 66.92555, 66.92294, 66.92034, 66.91772, 66.9151, 66.91249, 
    66.90989, 66.90726, 66.90462, 66.902, 66.89937, 66.89674, 66.89409, 
    66.89145, 66.88882, 66.88617, 66.88354, 66.88089, 66.87823, 66.87559, 
    66.87292,
  67.01666, 67.01414, 67.01159, 67.00905, 67.0065, 67.00396, 67.0014, 
    66.99884, 66.99628, 66.99373, 66.99115, 66.98859, 66.98603, 66.98344, 
    66.98088, 66.97829, 66.97571, 66.97312, 66.97053, 66.96793, 66.96531, 
    66.96272, 66.96012, 66.95751, 66.95491, 66.9523, 66.94968, 66.94706, 
    66.94445, 66.94183, 66.93921, 66.93656, 66.93394, 66.93131, 66.92867, 
    66.92604, 66.92342, 66.92076, 66.91811, 66.91547, 66.91281, 66.91015, 
    66.9075, 66.90485, 66.90219, 66.89954, 66.89687, 66.8942, 66.89153, 
    66.88885,
  67.0026, 67.0002, 66.9978, 66.99538, 66.99297, 66.99055, 66.98813, 
    66.98571, 66.98327, 66.98083, 66.9784, 66.97595, 66.9735, 66.97105, 
    66.9686, 66.96615, 66.96368, 66.96121, 66.95875, 66.95628, 66.95377, 
    66.95129, 66.94881, 66.94633, 66.94383, 66.94135, 66.93885, 66.93635, 
    66.93385, 66.93134, 66.92883, 66.92632, 66.92381, 66.92129, 66.91876, 
    66.91624, 66.91372, 66.91119, 66.90865, 66.90611, 66.90356, 66.90102, 
    66.89848, 66.89594, 66.89339, 66.89084, 66.88828, 66.88571, 66.88316, 
    66.88058,
  67.01941, 67.01699, 67.01456, 67.01212, 67.0097, 67.00726, 67.00482, 
    67.00238, 66.99992, 66.99746, 66.995, 66.99255, 66.99008, 66.98761, 
    66.98513, 66.98266, 66.98018, 66.9777, 66.97521, 66.97272, 66.9702, 
    66.9677, 66.96519, 66.9627, 66.96019, 66.95768, 66.95516, 66.95265, 
    66.95013, 66.94759, 66.94507, 66.94255, 66.94001, 66.93748, 66.93494, 
    66.9324, 66.92985, 66.92731, 66.92477, 66.92221, 66.91962, 66.91707, 
    66.91451, 66.91196, 66.90938, 66.90681, 66.90424, 66.90167, 66.89909, 
    66.89652,
  67.03622, 67.03377, 67.03133, 67.02888, 67.02643, 67.02397, 67.02151, 
    67.01904, 67.01656, 67.01408, 67.01161, 67.00914, 67.00665, 67.00417, 
    67.00166, 66.99918, 66.99667, 66.99418, 66.99166, 66.98916, 66.98663, 
    66.98411, 66.98159, 66.97906, 66.97653, 66.974, 66.97147, 66.96894, 
    66.96642, 66.96387, 66.96133, 66.95877, 66.95621, 66.95367, 66.9511, 
    66.94855, 66.94601, 66.94344, 66.94087, 66.9383, 66.9357, 66.93313, 
    66.93055, 66.92797, 66.92538, 66.9228, 66.9202, 66.91762, 66.91502, 
    66.91244,
  67.05302, 67.05056, 67.0481, 67.04563, 67.04316, 67.04068, 67.03819, 
    67.03571, 67.03322, 67.03072, 67.02823, 67.02573, 67.02322, 67.02072, 
    67.0182, 67.01569, 67.01318, 67.01066, 67.00813, 67.00561, 67.00307, 
    67.00052, 66.99798, 66.99543, 66.99288, 66.99033, 66.98779, 66.98524, 
    66.98269, 66.98013, 66.97757, 66.975, 66.97244, 66.96987, 66.96729, 
    66.96472, 66.96214, 66.95957, 66.95699, 66.95439, 66.95178, 66.94919, 
    66.94659, 66.94399, 66.94138, 66.93878, 66.93617, 66.93358, 66.93095, 
    66.92834,
  67.06982, 67.06735, 67.06487, 67.06238, 67.05988, 67.05738, 67.05489, 
    67.05238, 67.04987, 67.04736, 67.04484, 67.04231, 67.0398, 67.03728, 
    67.03474, 67.03221, 67.02967, 67.02713, 67.02459, 67.02203, 67.01949, 
    67.01694, 67.01437, 67.0118, 67.00925, 67.00668, 67.0041, 67.00155, 
    66.99897, 66.99639, 66.9938, 66.99123, 66.98865, 66.98606, 66.98347, 
    66.98088, 66.97829, 66.97568, 66.97308, 66.97044, 66.96785, 66.96523, 
    66.96262, 66.96002, 66.9574, 66.95477, 66.95214, 66.94953, 66.9469, 
    66.94427,
  67.08664, 67.08413, 67.08163, 67.07911, 67.07661, 67.07408, 67.07157, 
    67.06905, 67.06651, 67.06398, 67.06146, 67.05891, 67.05637, 67.05383, 
    67.05128, 67.04872, 67.04617, 67.04361, 67.04105, 67.03848, 67.03592, 
    67.03333, 67.03077, 67.02819, 67.0256, 67.02301, 67.02043, 67.01785, 
    67.01526, 67.01266, 67.01006, 67.00748, 67.00487, 67.00227, 66.99965, 
    66.99704, 66.99442, 66.99181, 66.98918, 66.98654, 66.9839, 66.98129, 
    66.97866, 66.97604, 66.9734, 66.97076, 66.96811, 66.96547, 66.96283, 
    66.96019,
  67.10343, 67.10093, 67.09839, 67.09586, 67.09334, 67.0908, 67.08826, 
    67.08571, 67.08316, 67.08061, 67.07806, 67.07551, 67.07294, 67.07039, 
    67.06781, 67.06524, 67.06267, 67.06009, 67.05752, 67.05492, 67.05235, 
    67.04974, 67.04716, 67.04457, 67.04196, 67.03937, 67.03677, 67.03416, 
    67.03155, 67.02892, 67.02631, 67.0237, 67.02106, 67.01845, 67.01583, 
    67.0132, 67.01056, 67.00793, 67.00529, 67.00265, 66.99999, 66.99734, 
    66.99471, 66.99204, 66.98938, 66.98674, 66.98408, 66.98142, 66.97876, 
    66.97612,
  67.12025, 67.11771, 67.11517, 67.11261, 67.11006, 67.10751, 67.10495, 
    67.10239, 67.09982, 67.09725, 67.09467, 67.09209, 67.08952, 67.08694, 
    67.08435, 67.08176, 67.07918, 67.07658, 67.07397, 67.07137, 67.06878, 
    67.06616, 67.06355, 67.06094, 67.05833, 67.05569, 67.05307, 67.05046, 
    67.04784, 67.04519, 67.04257, 67.03992, 67.03728, 67.03464, 67.032, 
    67.02935, 67.0267, 67.02405, 67.02141, 67.01874, 67.01608, 67.01343, 
    67.01076, 67.00809, 67.00542, 67.00274, 67.00006, 66.99738, 66.99471, 
    66.99203,
  67.10621, 67.1038, 67.10139, 67.09898, 67.09655, 67.09411, 67.09168, 
    67.08926, 67.08682, 67.08437, 67.08192, 67.07948, 67.07701, 67.07455, 
    67.0721, 67.06963, 67.06716, 67.06468, 67.06221, 67.05972, 67.05724, 
    67.05475, 67.05226, 67.04977, 67.04726, 67.04477, 67.04224, 67.03976, 
    67.03725, 67.03473, 67.0322, 67.02968, 67.02715, 67.02464, 67.0221, 
    67.01955, 67.01703, 67.01449, 67.01196, 67.0094, 67.00686, 67.00431, 
    67.00174, 66.99918, 66.99662, 66.99406, 66.99149, 66.98891, 66.98636, 
    66.98378,
  67.12302, 67.12059, 67.11815, 67.11572, 67.11327, 67.11083, 67.10838, 
    67.10593, 67.10346, 67.101, 67.09853, 67.09606, 67.09359, 67.09111, 
    67.08862, 67.08615, 67.08365, 67.08117, 67.07867, 67.07616, 67.07368, 
    67.07117, 67.06865, 67.06613, 67.06362, 67.0611, 67.05857, 67.05605, 
    67.05352, 67.05099, 67.04845, 67.0459, 67.04336, 67.04082, 67.03827, 
    67.03573, 67.03318, 67.03061, 67.02805, 67.02549, 67.02293, 67.02036, 
    67.01779, 67.01522, 67.01264, 67.01006, 67.00747, 67.00489, 67.0023, 
    66.99971 ;

 Longitude =
  46.51716, 46.47765, 46.43822, 46.39891, 46.35968, 46.32058, 46.28156, 
    46.24268, 46.20383, 46.16513, 46.12648, 46.08799, 46.04957, 46.01125, 
    45.97302, 45.93488, 45.89684, 45.85889, 45.82104, 45.78316, 45.74537, 
    45.70775, 45.67018, 45.63273, 45.59543, 45.55842, 45.52107, 45.48421, 
    45.44712, 45.41035, 45.37339, 45.33672, 45.30018, 45.26367, 45.22721, 
    45.19092, 45.15468, 45.11847, 45.08233, 45.0463, 45.0104, 44.97458, 
    44.93879, 44.90312, 44.86756, 44.83205, 44.7967, 44.76129, 44.72601, 
    44.69084,
  46.51044, 46.47093, 46.43146, 46.39213, 46.35291, 46.31378, 46.27477, 
    46.23582, 46.19698, 46.15827, 46.1196, 46.08109, 46.04266, 46.00429, 
    45.96606, 45.92792, 45.88983, 45.85188, 45.81401, 45.77608, 45.73838, 
    45.70064, 45.66307, 45.6256, 45.58849, 45.55126, 45.51389, 45.47682, 
    45.43988, 45.40301, 45.36617, 45.32946, 45.29288, 45.25637, 45.21996, 
    45.18361, 45.14734, 45.11115, 45.07497, 45.03897, 45.00304, 44.96717, 
    44.93139, 44.89571, 44.86007, 44.82462, 44.78921, 44.75384, 44.71856, 
    44.68334,
  46.50376, 46.4642, 46.42477, 46.3854, 46.34613, 46.30702, 46.26795, 
    46.22897, 46.19012, 46.15139, 46.11274, 46.07417, 46.03571, 45.99737, 
    45.95909, 45.92092, 45.88286, 45.84486, 45.80696, 45.76916, 45.73118, 
    45.69353, 45.656, 45.61853, 45.58119, 45.54401, 45.50673, 45.46965, 
    45.4327, 45.39584, 45.35898, 45.32223, 45.28561, 45.2491, 45.21268, 
    45.17628, 45.14002, 45.10387, 45.0677, 45.03166, 44.99564, 44.95973, 
    44.92397, 44.88835, 44.85266, 44.81717, 44.78171, 44.74647, 44.71105, 
    44.67587,
  46.49706, 46.4575, 46.41802, 46.37867, 46.33934, 46.3002, 46.26112, 
    46.22216, 46.18331, 46.14454, 46.10584, 46.06729, 46.02881, 45.99043, 
    45.95215, 45.91393, 45.87587, 45.83783, 45.79993, 45.76213, 45.72405, 
    45.68644, 45.64888, 45.6114, 45.57404, 45.5368, 45.49961, 45.46247, 
    45.42551, 45.38857, 45.35173, 45.315, 45.27835, 45.24184, 45.2054, 
    45.16902, 45.1327, 45.09652, 45.06042, 45.02434, 44.98829, 44.95233, 
    44.91651, 44.88089, 44.84529, 44.80976, 44.77428, 44.73893, 44.70355, 
    44.66837,
  46.49037, 46.45079, 46.41129, 46.37187, 46.3326, 46.2934, 46.25431, 
    46.21533, 46.17643, 46.13766, 46.09896, 46.06038, 46.0219, 45.98349, 
    45.94519, 45.90698, 45.86888, 45.83084, 45.79289, 45.75507, 45.71702, 
    45.6793, 45.64178, 45.60431, 45.56693, 45.52969, 45.49246, 45.45532, 
    45.41832, 45.38138, 45.34452, 45.30773, 45.27111, 45.23458, 45.19812, 
    45.16173, 45.12548, 45.08923, 45.05308, 45.01699, 44.98087, 44.94493, 
    44.90912, 44.87342, 44.83788, 44.80236, 44.76681, 44.73148, 44.69611, 
    44.66084,
  46.48796, 46.44836, 46.40884, 46.36943, 46.33012, 46.29089, 46.25177, 
    46.21277, 46.17385, 46.135, 46.09629, 46.05765, 46.0191, 45.98069, 
    45.94237, 45.90414, 45.86597, 45.8279, 45.78996, 45.75208, 45.71393, 
    45.67624, 45.63869, 45.60113, 45.56373, 45.52641, 45.48923, 45.45203, 
    45.41501, 45.37803, 45.34114, 45.30436, 45.26765, 45.23102, 45.19456, 
    45.15812, 45.1218, 45.08555, 45.04933, 45.01323, 44.97704, 44.94106, 
    44.90522, 44.86953, 44.8339, 44.79831, 44.76278, 44.72733, 44.69194, 
    44.65674,
  46.48121, 46.44161, 46.40201, 46.36259, 46.32327, 46.28403, 46.24491, 
    46.20587, 46.16694, 46.1281, 46.08931, 46.0507, 46.01215, 45.97369, 
    45.93533, 45.8971, 45.85892, 45.82085, 45.78287, 45.74502, 45.70689, 
    45.66911, 45.63155, 45.59402, 45.55653, 45.51917, 45.48196, 45.44482, 
    45.40776, 45.37074, 45.33387, 45.29706, 45.26037, 45.22378, 45.18723, 
    45.15082, 45.11447, 45.07821, 45.04203, 45.00587, 44.9696, 44.93362, 
    44.89776, 44.862, 44.82638, 44.79074, 44.7552, 44.71975, 44.68435, 
    44.64914,
  46.47445, 46.43481, 46.39523, 46.35578, 46.31645, 46.27718, 46.23805, 
    46.19898, 46.16003, 46.12115, 46.0824, 46.04374, 46.00518, 45.96668, 
    45.92833, 45.89005, 45.85187, 45.81379, 45.77577, 45.73788, 45.7, 
    45.66203, 45.62439, 45.58674, 45.54924, 45.51189, 45.47466, 45.43754, 
    45.4005, 45.36353, 45.32663, 45.28977, 45.25304, 45.21648, 45.17994, 
    45.14348, 45.10715, 45.07089, 45.03468, 44.99853, 44.96211, 44.92618, 
    44.89035, 44.85452, 44.81884, 44.78321, 44.74763, 44.71222, 44.67678, 
    44.64156,
  46.46774, 46.42803, 46.38847, 46.349, 46.30959, 46.27036, 46.23119, 
    46.1921, 46.15311, 46.11423, 46.07547, 46.03678, 45.99818, 45.95971, 
    45.92131, 45.88303, 45.84484, 45.80672, 45.7687, 45.7308, 45.69297, 
    45.65496, 45.61721, 45.57953, 45.54199, 45.50467, 45.4674, 45.43033, 
    45.39324, 45.35626, 45.31938, 45.28255, 45.24584, 45.20921, 45.17266, 
    45.13616, 45.09975, 45.06353, 45.02736, 44.99102, 44.95473, 44.91871, 
    44.88289, 44.84711, 44.81134, 44.77565, 44.74007, 44.70466, 44.66924, 
    44.63398,
  46.46096, 46.42129, 46.38168, 46.34217, 46.3028, 46.26353, 46.2243, 
    46.18523, 46.14624, 46.10734, 46.06855, 46.0298, 45.99124, 45.95272, 
    45.91432, 45.876, 45.83778, 45.79965, 45.76162, 45.72369, 45.68584, 
    45.64791, 45.61023, 45.57264, 45.53516, 45.49773, 45.46037, 45.42318, 
    45.38606, 45.34904, 45.31212, 45.27531, 45.23858, 45.20193, 45.16534, 
    45.12879, 45.09252, 45.05608, 45.01977, 44.98337, 44.94724, 44.91127, 
    44.87539, 44.8396, 44.80383, 44.76819, 44.73257, 44.69706, 44.66162, 
    44.62637,
  46.45421, 46.41452, 46.37491, 46.33535, 46.29597, 46.25666, 46.21746, 
    46.17834, 46.13935, 46.10041, 46.0616, 46.02287, 45.98426, 45.94574, 
    45.90729, 45.86897, 45.83074, 45.79258, 45.75454, 45.71657, 45.67871, 
    45.64074, 45.60308, 45.56553, 45.52799, 45.49059, 45.45332, 45.41608, 
    45.37896, 45.34194, 45.30492, 45.26806, 45.23124, 45.19455, 45.15796, 
    45.12145, 45.0851, 45.04873, 45.01234, 44.97583, 44.93963, 44.9036, 
    44.86778, 44.83204, 44.79626, 44.76054, 44.72491, 44.68941, 44.65396, 
    44.61865,
  46.44748, 46.40775, 46.36811, 46.32855, 46.28916, 46.24984, 46.21058, 
    46.17145, 46.1324, 46.09347, 46.05466, 46.0159, 45.97726, 45.93874, 
    45.90028, 45.86193, 45.82369, 45.78552, 45.74743, 45.70947, 45.67162, 
    45.63373, 45.59599, 45.55838, 45.52083, 45.48341, 45.4461, 45.40893, 
    45.37176, 45.33461, 45.29758, 45.26074, 45.22393, 45.18722, 45.15061, 
    45.11406, 45.07758, 45.04121, 45.00496, 44.96866, 44.93242, 44.89632, 
    44.86033, 44.82442, 44.78865, 44.75291, 44.71729, 44.68173, 44.6463, 
    44.61107,
  46.44075, 46.40099, 46.36134, 46.32178, 46.28231, 46.24298, 46.20371, 
    46.16458, 46.12554, 46.0866, 46.04771, 46.00896, 45.97029, 45.93174, 
    45.89328, 45.8549, 45.81663, 45.77845, 45.74034, 45.70236, 45.66445, 
    45.62667, 45.58892, 45.55122, 45.51371, 45.47617, 45.43881, 45.40163, 
    45.3645, 45.32739, 45.2904, 45.2534, 45.21656, 45.17982, 45.14317, 
    45.10662, 45.07013, 45.03378, 44.9975, 44.96126, 44.92519, 44.8891, 
    44.85311, 44.81726, 44.78141, 44.74559, 44.70991, 44.67424, 44.63876, 
    44.60345,
  46.43872, 46.39893, 46.35923, 46.31966, 46.28017, 46.24077, 46.2015, 
    46.16228, 46.12324, 46.08423, 46.04535, 46.00655, 45.96787, 45.92928, 
    45.89077, 45.85236, 45.81405, 45.77584, 45.73773, 45.69971, 45.66179, 
    45.62389, 45.5861, 45.54845, 45.51088, 45.47339, 45.43597, 45.39874, 
    45.36154, 45.32435, 45.28721, 45.25024, 45.21344, 45.17671, 45.14, 
    45.10344, 45.06689, 45.03051, 44.99417, 44.9579, 44.92175, 44.88565, 
    44.84954, 44.81355, 44.77764, 44.74189, 44.70619, 44.67055, 44.63511, 
    44.5997,
  46.4319, 46.39211, 46.35241, 46.31281, 46.2733, 46.23388, 46.19458, 
    46.1554, 46.11628, 46.07727, 46.03837, 45.99955, 45.96085, 45.92221, 
    45.88371, 45.84529, 45.80696, 45.76873, 45.73058, 45.69256, 45.65462, 
    45.61675, 45.5789, 45.54121, 45.50367, 45.46609, 45.4286, 45.39139, 
    45.35415, 45.31709, 45.27998, 45.243, 45.20608, 45.16926, 45.13259, 
    45.09597, 45.05947, 45.02301, 44.98663, 44.95044, 44.9143, 44.8782, 
    44.84216, 44.80625, 44.77032, 44.73455, 44.69887, 44.66325, 44.62769, 
    44.59214 ;

 MaxIceConc = 100 ;

 MeanIceConc = 88.47009 ;

 MinIceConc = 14.89622 ;

 NumOfQACategories = 4 ;

 QCFlags =
  -20905760, -20905760, -20905760, -20905760, -17760030, -20905760, 
    -20905751, -20905751, -20905751, -16973662, -16973662, -16973594, 
    -17497878, -16973662, -16973594, -16973594, -16973594, -16908058, 
    -16908062, -16908054, -16908054, -16908054, -16908054, -16908054, 
    -16908062, -16908054, -16908054, -16908054, -17301270, -16908054, 
    -16908054, -16908054, -16908062, -16908054, -16908054, -16908054, 
    -16908054, -16908054, -16908058, -16908058, -16908050, -16908050, 
    -16908050, -16908050, -16908050, -16908050, -16908050, -16908050, 
    -16908050, -16908050,
  -20905751, -20905751, -20905751, -17760030, -20905760, -20905760, 
    -20905760, -20905760, -20905760, -20905760, -20905751, -16973662, 
    -16973594, -17760030, -16973662, -16973594, -17497878, -16908058, 
    -16908058, -16908054, -16908054, -16908054, -16908054, -16908054, 
    -16908054, -16908054, -16908054, -16908054, -16908054, -16908054, 
    -16908054, -16908054, -16908062, -16908054, -16908054, -16908054, 
    -16908054, -16908054, -16908054, -16908054, -16908058, -16908058, 
    -16908058, -16908058, -16908050, -16908050, -16908050, -16908050, 
    -16908050, -16908050,
  -17760022, -16973594, -17760022, -20905751, -20905760, -16973594, 
    -20905760, -20905760, -20905760, -20905760, -20905760, -20905760, 
    -17760022, -17760022, -16973662, -16973594, -17497878, -16908058, 
    -16908058, -16908058, -16908054, -16908054, -16908054, -16908054, 
    -16908054, -16908054, -16908054, -16908054, -16908054, -16908054, 
    -16908054, -16908062, -16908062, -16908054, -16908054, -16908054, 
    -16908054, -16908054, -16908054, -16908054, -16908054, -16908054, 
    -16908054, -16908054, -16908126, -16908050, -16908050, -16908050, 
    -16908050, -16908050,
  -16973594, -16973586, -16973594, -16973594, -20905751, -16973662, 
    -17760030, -17760030, -17760030, -20905751, -20905760, -16973662, 
    -20905760, -17760022, -17760030, -16973594, -16973594, -16973594, 
    -16908058, -16908058, -16908054, -16908054, -16908054, -16908054, 
    -16908054, -16908054, -16908054, -16908054, -16908054, -16908054, 
    -16908054, -16908062, -16908062, -16908054, -16908054, -16908054, 
    -16908054, -16908054, -16908054, -16908054, -16908054, -16908054, 
    -16908054, -16908054, -16908126, -16908126, -16908058, -16908050, 
    -16908050, -16908050,
  -16973586, -17760022, -17760022, -16973594, -20905760, -20905751, 
    -17760030, -20905760, -17760030, -20905760, -20905760, -20905760, 
    -16973662, -17760030, -17760030, -17497886, -16973662, -16973662, 
    -17497886, -16908062, -16908054, -16908054, -16908054, -16908054, 
    -16908054, -16908054, -16908054, -16908054, -16908054, -16908054, 
    -16908054, -16908062, -16908062, -16908062, -16908054, -16908054, 
    -16908054, -16908054, -16908054, -16908054, -16908054, -16908054, 
    -16908054, -16908062, -16908126, -16908126, -16908054, -16908054, 
    -16908050, -16908050,
  -16973594, -16973594, -16973594, -20905751, -20905751, -20905751, 
    -17760022, -20905760, -17497886, -20905760, -20905760, -20905760, 
    -16973662, -17760030, -17760022, -17497886, -16973594, -16973594, 
    -16908126, -16908126, -16908054, -16908054, -16908054, -16908054, 
    -16908054, -16908054, -16908054, -16908054, -16908054, -16908054, 
    -16908054, -16908062, -16908062, -16908054, -16908054, -16908054, 
    -16908054, -16908054, -16908054, -16908054, -16908054, -16908054, 
    -16908054, -16908062, -16908062, -16908062, -16908050, -16908126, 
    -16908050, -16908050,
  -20905751, -16973594, -16973594, -16973594, -20905751, -20905751, 
    -20905760, -20905751, -17760030, -20905751, -20905751, -20905751, 
    -20905751, -17760030, -20905760, -17760030, -16973594, -16973594, 
    -16908058, -16908062, -16908054, -16908054, -16908054, -16908054, 
    -16908054, -16908054, -16908054, -16908054, -16908054, -16908054, 
    -16908054, -16908062, -16908062, -16908054, -16908054, -16908054, 
    -16908054, -16908054, -16908054, -16908058, -16908054, -16908062, 
    -16908062, -16908062, -16908050, -16908062, -16908126, -16908126, 
    -16908050, -16908050,
  -16973662, -20905751, -20905751, -16973662, -16973594, -20905751, 
    -17760022, -20905751, -17760030, -20905751, -17760030, -20905751, 
    -20905751, -20905751, -20905751, -20905760, -20905760, -17760030, 
    -16973662, -16908058, -16908054, -16908054, -16908054, -16908054, 
    -16908062, -16908054, -16908054, -16908054, -16908054, -16908054, 
    -16908062, -16908062, -16908062, -16908054, -16908054, -16908054, 
    -16908054, -16908054, -16908054, -16908054, -16908058, -16908054, 
    -16908054, -16908054, -16908050, -16908058, -16908050, -16908050, 
    -16908058, -16908058,
  -20905760, -20905760, -20905760, -20905760, -16973662, -16973594, 
    -20905751, -20905760, -20905751, -20905760, -17760030, -17760030, 
    -20905760, -20905760, -20905751, -20905751, -20905760, -20905760, 
    -20905760, -16973594, -16908058, -16908054, -16908054, -16908054, 
    -16908054, -16908054, -16908054, -16908054, -16908062, -16908062, 
    -16908062, -16908062, -16908062, -16908054, -16908054, -16908054, 
    -16908054, -16908054, -16908054, -16908054, -16908054, -16908054, 
    -16908054, -16908050, -16908054, -16908054, -16908054, -16908050, 
    -16908058, -16908054,
  -20905760, -20905760, -20905760, -20905760, -20905760, -16973662, 
    -20905751, -20905751, -16973586, -16973586, -17497878, -17760022, 
    -17760030, -20905760, -20905760, -20905760, -20905760, -20905760, 
    -17760030, -16908126, -16908058, -16908054, -16908054, -16908054, 
    -16908054, -16908054, -16908054, -16908054, -16908054, -16908054, 
    -16908054, -16908062, -16908062, -16908054, -16908054, -16908054, 
    -17039126, -16908054, -16908054, -16908054, -16908054, -16908054, 
    -16908054, -16908050, -16908050, -16908054, -16908054, -16908054, 
    -16908062, -16908054,
  -20905760, -20905760, -20905760, -20905760, -20905760, -20905760, 
    -20905760, -16973662, -20905751, -20905760, -17497878, -16973586, 
    -20905760, -20905760, -20905760, -20905760, -17760030, -20905760, 
    -17497886, -16908062, -16908058, -16908054, -16908054, -16908054, 
    -16908054, -16908054, -16908054, -16908054, -16908054, -16908054, 
    -16908054, -16908062, -16908054, -16908054, -16908054, -16908054, 
    -16908054, -16908054, -16908054, -16908054, -16908054, -16908054, 
    -16908054, -16908054, -16908058, -16908054, -16908058, -16908058, 
    -16908054, -16908054,
  -20905760, -20905760, -20905760, -20905760, -20905760, -20905760, 
    -20905760, -16973662, -16973662, -20905760, -16973662, -20905760, 
    -17497886, -17497886, -20905760, -20905760, -20905760, -17497886, 
    -16973594, -16973594, -16908062, -16908054, -16908054, -16908054, 
    -16908054, -16908054, -16908054, -16908054, -16908054, -16908054, 
    -16908054, -16908054, -16908054, -16908054, -16908054, -16908054, 
    -16908054, -16908054, -16908054, -16908054, -16908054, -16908054, 
    -16908054, -16908054, -16908054, -16908054, -16908054, -16908054, 
    -16908050, -16908050,
  -20905760, -20905760, -20905760, -20905760, -20905760, -16973586, 
    -16973662, -20905760, -20905760, -20905760, -20905760, -20905760, 
    -20905760, -16973586, -16973586, -18546454, -16973662, -18546462, 
    -18546462, -17497886, -16908062, -16908054, -16908054, -16908054, 
    -16908054, -16908054, -16908054, -16908054, -16908054, -16908054, 
    -16908054, -16908054, -16908054, -16908054, -16908054, -16908054, 
    -16908054, -16908054, -16908054, -17301270, -16908062, -16908062, 
    -16908054, -16908054, -16908054, -16908054, -16908054, -16908126, 
    -16908050, -16908050,
  -20905760, -20905760, -20905760, -20905760, -20905760, -16973594, 
    -20905760, -20905760, -20905760, -20905760, -20905760, -20905760, 
    -20905751, -17497878, -16973594, -18546462, -16973662, -17497886, 
    -18546462, -16908062, -16908062, -16908054, -16908054, -16908054, 
    -16908054, -16908054, -16908054, -16908054, -16908054, -16908054, 
    -16908054, -16908054, -16908054, -16908054, -16908054, -16908054, 
    -16908054, -16908054, -16908054, -16908054, -16908062, -16908062, 
    -16908054, -16908054, -16908054, -16908054, -16908054, -16908126, 
    -16908050, -16908058,
  -20905760, -20905760, -20905760, -20905760, -20905760, -20905751, 
    -20905760, -20905760, -20905760, -20905760, -20905760, -18546462, 
    -20905760, -16973586, -16973586, -16973594, -16973662, -17497886, 
    -18546462, -17497886, -16908062, -16908054, -16908054, -16908054, 
    -16908054, -16908054, -16908054, -16908054, -16908054, -16908054, 
    -16908054, -16908054, -16908054, -16908054, -16908054, -16908054, 
    -16908054, -16908054, -16908054, -17301270, -17301270, -16908054, 
    -17039126, -16908054, -16908054, -16908054, -16908054, -16908062, 
    -16908054, -16908054 ;

 STDIceConc = 19.20647 ;

 SearchWindowSize = 50 ;

 StartColumn = 1 ;

 StartRow = 1 ;

 SummaryQC_Ice_Concentration =
  0, 0, 0, 0, 2, 0, 1, 1, 1, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  1, 1, 1, 2, 0, 0, 0, 0, 0, 0, 1, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  2, 2, 2, 1, 0, 2, 0, 0, 0, 0, 0, 0, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  2, 2, 2, 2, 1, 2, 2, 2, 2, 1, 0, 2, 0, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  2, 2, 2, 2, 0, 1, 2, 0, 2, 0, 0, 0, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  2, 2, 2, 1, 1, 1, 2, 0, 2, 0, 0, 0, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  1, 2, 2, 2, 1, 1, 0, 1, 2, 1, 1, 1, 1, 2, 0, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  2, 1, 1, 2, 2, 1, 2, 1, 2, 1, 2, 1, 1, 1, 1, 0, 0, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  0, 0, 0, 0, 2, 2, 1, 0, 1, 0, 2, 2, 0, 0, 1, 1, 0, 0, 0, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  0, 0, 0, 0, 0, 2, 1, 1, 2, 2, 2, 2, 2, 0, 0, 0, 0, 0, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  0, 0, 0, 0, 0, 0, 0, 2, 1, 0, 2, 2, 0, 0, 0, 0, 2, 0, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  0, 0, 0, 0, 0, 0, 0, 2, 2, 0, 2, 0, 2, 2, 0, 0, 0, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  0, 0, 0, 0, 0, 2, 2, 0, 0, 0, 0, 0, 0, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 1, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 2, 0, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2 ;

 TotDaytimePixs = 6731 ;

 TotIceRetrvls = 6731 ;

 TotIceTermnt = 2450869 ;

 TotNighttimePixs = _ ;

 TotWaterPixs = 114350 ;

 Tot_QA_BadData = 55710 ;

 Tot_QA_Nonretrievable = 2395159 ;

 Tot_QA_Normal = 5596 ;

 Tot_QA_Uncertain = 1135 ;
}
