netcdf sss_smos_2_sub {
dimensions:
	n_grid_points = 52 ;
variables:
	short Dg_quality_SSS_corr(n_grid_points) ;
		Dg_quality_SSS_corr:_FillValue = 999US ;
		string Dg_quality_SSS_corr:_Unsigned = "true" ;
	float Latitude(n_grid_points) ;
		string Latitude:units = "deg" ;
		Latitude:_FillValue = -999.f ;
	float Longitude(n_grid_points) ;
		string Longitude:units = "deg" ;
		Longitude:_FillValue = -999.f ;
	float Mean_acq_time(n_grid_points) ;
		string Mean_acq_time:units = "dd" ;
		Mean_acq_time:_FillValue = -999.f ;
	float SSS_corr(n_grid_points) ;
		string SSS_corr:units = "psu" ;
		SSS_corr:_FillValue = -999.f ;
	float Sigma_SSS_corr(n_grid_points) ;
		string Sigma_SSS_corr:units = "psu" ;
		Sigma_SSS_corr:_FillValue = -999.f ;

// global attributes:
		string :creation_date = "UTC=2021-07-01T05:16:26" ;
		string :total_number_of_grid_points = "92713" ;
		string :FH\:File_Name = "SM_OPER_MIR_OSUDP2_20210630T215911_20210630T225230_700_001_1" ;
		string :FH\:File_Description = "L2 Ocean Salinity Output User Data Product." ;
		string :FH\:Notes = "The UDP (User Data Product) is designed for oceanographics and high level centers, it includes geophysical parameters, a theoretical estimate of their accuracy, flags and descriptors of the product quality." ;
		string :FH\:Mission = "SMOS" ;
		string :FH\:File_Class = "OPER" ;
		string :FH\:File_Type = "MIR_OSUDP2" ;
		string :FH\:File_Version = "0001" ;
		string :FH\:Validity_Period\:Validity_Start = "UTC=2021-06-30T21:59:11" ;
		string :FH\:Validity_Period\:Validity_Stop = "UTC=2021-06-30T22:52:30" ;
		string :FH\:Source\:System = "DPGS" ;
		string :FH\:Source\:Creator = "L2OP" ;
		string :FH\:Source\:Creator_Version = "700" ;
		string :FH\:Source\:Creation_Date = "UTC=2021-07-01T05:09:30" ;
		string :VH\:SPH\:QI\:Total_Selected_L1c_Grid_Points = "60219" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:Retrieval_Scheme = "1" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:Land_Rejected = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:Too_Close_To_Land_Rejected = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:Ice_Rejected = "10855" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:Missing_ECMWF_Rejected = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:Too_Few_Measurements_Rejected = "18084" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:Good_Quality_Grid_Points = "29636" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:Poor_Quality_Grid_Points = "4896" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:SQ\:Grid_Point_Type = "Sea" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:SQ\:SSS_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:SQ\:SST_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:SQ\:WS_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:SQ\:Good_Quality = "23293" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:SQ\:Good_Quality_Retrieved = "17816" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:SQ\:Good_Quality_Retrieved_Average_Sigma = "1.959542" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:SQ\:Good_Quality_Failed_Outside_Valid_Range = "81" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:SQ\:Good_Quality_Failed_Sigma_Too_High = "478" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:SQ\:Good_Quality_Failed_Poor_Fit = "5037" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:SQ\:Good_Quality_Failed_Marquardt = "4" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:SQ\:Good_Quality_Failed_Maxiter = "110" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:SQ\:Good_Quality_Failed_OOLUT = "555" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:SQ\:Poor_Quality = "2426" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:SQ\:Poor_Quality_Retrieved = "1661" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:SQ\:Poor_Quality_Retrieved_Average_Sigma = "2.933723" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:NCQ\:Grid_Point_Type = "Near_Coast" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:NCQ\:SSS_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:NCQ\:SST_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:NCQ\:WS_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:NCQ\:Good_Quality = "6343" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:NCQ\:Good_Quality_Retrieved = "3803" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:NCQ\:Good_Quality_Retrieved_Average_Sigma = "1.253443" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:NCQ\:Good_Quality_Failed_Outside_Valid_Range = "276" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:NCQ\:Good_Quality_Failed_Sigma_Too_High = "522" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:NCQ\:Good_Quality_Failed_Poor_Fit = "2247" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:NCQ\:Good_Quality_Failed_Marquardt = "152" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:NCQ\:Good_Quality_Failed_Maxiter = "411" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:NCQ\:Good_Quality_Failed_OOLUT = "773" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:NCQ\:Poor_Quality = "2470" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:NCQ\:Poor_Quality_Retrieved = "1367" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:NCQ\:Poor_Quality_Retrieved_Average_Sigma = "1.480500" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_0\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_0\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_0\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_0\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_0\:Good_Quality = "559" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_0\:Good_Quality_Retrieved = "131" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_0\:Good_Quality_Retrieved_Average_Sigma = "1.985529" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_0\:Good_Quality_Failed_Outside_Valid_Range = "183" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_0\:Good_Quality_Failed_Sigma_Too_High = "261" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_0\:Good_Quality_Failed_Poor_Fit = "325" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_0\:Good_Quality_Failed_Marquardt = "112" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_0\:Good_Quality_Failed_Maxiter = "130" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_0\:Good_Quality_Failed_OOLUT = "326" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_0\:Poor_Quality = "106" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_0\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_0\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_1\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_1\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_1\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_1\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_1\:Good_Quality = "486" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_1\:Good_Quality_Retrieved = "229" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_1\:Good_Quality_Retrieved_Average_Sigma = "2.167454" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_1\:Good_Quality_Failed_Outside_Valid_Range = "60" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_1\:Good_Quality_Failed_Sigma_Too_High = "82" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_1\:Good_Quality_Failed_Poor_Fit = "244" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_1\:Good_Quality_Failed_Marquardt = "30" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_1\:Good_Quality_Failed_Maxiter = "45" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_1\:Good_Quality_Failed_OOLUT = "135" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_1\:Poor_Quality = "233" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_1\:Poor_Quality_Retrieved = "13" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_1\:Poor_Quality_Retrieved_Average_Sigma = "4.597799" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_2\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_2\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_2\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_2\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_2\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_2\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_2\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_2\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_2\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_2\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_2\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_2\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_2\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_2\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_2\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_2\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_3\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_3\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_3\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_3\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_3\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_3\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_3\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_3\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_3\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_3\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_3\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_3\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_3\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_3\:Poor_Quality = "3" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_3\:Poor_Quality_Retrieved = "1" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_3\:Poor_Quality_Retrieved_Average_Sigma = "2.726585" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_4\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_4\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_4\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_4\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_4\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_4\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_4\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_4\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_4\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_4\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_4\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_4\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_4\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_4\:Poor_Quality = "233" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_4\:Poor_Quality_Retrieved = "182" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_4\:Poor_Quality_Retrieved_Average_Sigma = "3.945308" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_5\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_5\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_5\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_5\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_5\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_5\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_5\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_5\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_5\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_5\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_5\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_5\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_5\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_5\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_5\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_5\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_6\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_6\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_6\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_6\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_6\:Good_Quality = "16" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_6\:Good_Quality_Retrieved = "14" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_6\:Good_Quality_Retrieved_Average_Sigma = "1.307737" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_6\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_6\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_6\:Good_Quality_Failed_Poor_Fit = "2" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_6\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_6\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_6\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_6\:Poor_Quality = "22" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_6\:Poor_Quality_Retrieved = "19" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_6\:Poor_Quality_Retrieved_Average_Sigma = "1.902701" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_7\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_7\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_7\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_7\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_7\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_7\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_7\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_7\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_7\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_7\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_7\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_7\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_7\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_7\:Poor_Quality = "113" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_7\:Poor_Quality_Retrieved = "58" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_7\:Poor_Quality_Retrieved_Average_Sigma = "1.925949" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_8\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_8\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_8\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_8\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_8\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_8\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_8\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_8\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_8\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_8\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_8\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_8\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_8\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_8\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_8\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_8\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_9\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_9\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_9\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_9\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_9\:Good_Quality = "1485" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_9\:Good_Quality_Retrieved = "825" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_9\:Good_Quality_Retrieved_Average_Sigma = "2.191673" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_9\:Good_Quality_Failed_Outside_Valid_Range = "1" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_9\:Good_Quality_Failed_Sigma_Too_High = "54" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_9\:Good_Quality_Failed_Poor_Fit = "544" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_9\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_9\:Good_Quality_Failed_Maxiter = "247" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_9\:Good_Quality_Failed_OOLUT = "190" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_9\:Poor_Quality = "11" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_9\:Poor_Quality_Retrieved = "1" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_9\:Poor_Quality_Retrieved_Average_Sigma = "4.534814" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_10\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_10\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_10\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_10\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_10\:Good_Quality = "6940" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_10\:Good_Quality_Retrieved = "4685" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_10\:Good_Quality_Retrieved_Average_Sigma = "2.611991" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_10\:Good_Quality_Failed_Outside_Valid_Range = "102" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_10\:Good_Quality_Failed_Sigma_Too_High = "600" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_10\:Good_Quality_Failed_Poor_Fit = "1779" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_10\:Good_Quality_Failed_Marquardt = "14" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_10\:Good_Quality_Failed_Maxiter = "72" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_10\:Good_Quality_Failed_OOLUT = "603" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_10\:Poor_Quality = "508" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_10\:Poor_Quality_Retrieved = "218" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_10\:Poor_Quality_Retrieved_Average_Sigma = "4.334874" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_11\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_11\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_11\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_11\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_11\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_11\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_11\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_11\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_11\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_11\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_11\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_11\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_11\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_11\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_11\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_11\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_12\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_12\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_12\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_12\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_12\:Good_Quality = "232" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_12\:Good_Quality_Retrieved = "156" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_12\:Good_Quality_Retrieved_Average_Sigma = "1.521774" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_12\:Good_Quality_Failed_Outside_Valid_Range = "1" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_12\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_12\:Good_Quality_Failed_Poor_Fit = "70" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_12\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_12\:Good_Quality_Failed_Maxiter = "7" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_12\:Good_Quality_Failed_OOLUT = "17" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_12\:Poor_Quality = "55" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_12\:Poor_Quality_Retrieved = "42" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_12\:Poor_Quality_Retrieved_Average_Sigma = "2.482193" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_13\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_13\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_13\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_13\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_13\:Good_Quality = "11990" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_13\:Good_Quality_Retrieved = "9532" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_13\:Good_Quality_Retrieved_Average_Sigma = "2.064730" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_13\:Good_Quality_Failed_Outside_Valid_Range = "10" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_13\:Good_Quality_Failed_Sigma_Too_High = "3" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_13\:Good_Quality_Failed_Poor_Fit = "2454" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_13\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_13\:Good_Quality_Failed_Maxiter = "1" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_13\:Good_Quality_Failed_OOLUT = "42" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_13\:Poor_Quality = "997" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_13\:Poor_Quality_Retrieved = "857" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_13\:Poor_Quality_Retrieved_Average_Sigma = "3.092174" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_14\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_14\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_14\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_14\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_14\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_14\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_14\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_14\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_14\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_14\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_14\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_14\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_14\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_14\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_14\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_14\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_15\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_15\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_15\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_15\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_15\:Good_Quality = "830" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_15\:Good_Quality_Retrieved = "677" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_15\:Good_Quality_Retrieved_Average_Sigma = "1.047869" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_15\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_15\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_15\:Good_Quality_Failed_Poor_Fit = "153" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_15\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_15\:Good_Quality_Failed_Maxiter = "1" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_15\:Good_Quality_Failed_OOLUT = "4" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_15\:Poor_Quality = "1379" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_15\:Poor_Quality_Retrieved = "1092" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_15\:Poor_Quality_Retrieved_Average_Sigma = "1.087475" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_16\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_16\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_16\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_16\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_16\:Good_Quality = "7097" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_16\:Good_Quality_Retrieved = "5369" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_16\:Good_Quality_Retrieved_Average_Sigma = "0.787403" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_16\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_16\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_16\:Good_Quality_Failed_Poor_Fit = "1713" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_16\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_16\:Good_Quality_Failed_Maxiter = "18" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_16\:Good_Quality_Failed_OOLUT = "11" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_16\:Poor_Quality = "1043" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_16\:Poor_Quality_Retrieved = "450" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_16\:Poor_Quality_Retrieved_Average_Sigma = "1.581808" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_17\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_17\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_17\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_17\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_17\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_17\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_17\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_17\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_17\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_17\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_17\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_17\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_17\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_17\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_17\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_17\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_18\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_18\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_18\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_18\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_18\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_18\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_18\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_18\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_18\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_18\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_18\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_18\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_18\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_18\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_18\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_18\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_19\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_19\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_19\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_19\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_19\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_19\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_19\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_19\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_19\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_19\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_19\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_19\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_19\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_19\:Poor_Quality = "141" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_19\:Poor_Quality_Retrieved = "51" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_19\:Poor_Quality_Retrieved_Average_Sigma = "4.372903" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_20\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_20\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_20\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_20\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_20\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_20\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_20\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_20\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_20\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_20\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_20\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_20\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_20\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_20\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_20\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_20\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_21\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_21\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_21\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_21\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_21\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_21\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_21\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_21\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_21\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_21\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_21\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_21\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_21\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_21\:Poor_Quality = "8" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_21\:Poor_Quality_Retrieved = "5" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_21\:Poor_Quality_Retrieved_Average_Sigma = "2.769263" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_22\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_22\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_22\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_22\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_22\:Good_Quality = "1" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_22\:Good_Quality_Retrieved = "1" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_22\:Good_Quality_Retrieved_Average_Sigma = "2.597888" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_22\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_22\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_22\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_22\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_22\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_22\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_22\:Poor_Quality = "42" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_22\:Poor_Quality_Retrieved = "37" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_22\:Poor_Quality_Retrieved_Average_Sigma = "3.355307" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_23\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_23\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_23\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_23\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_23\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_23\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_23\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_23\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_23\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_23\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_23\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_23\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_23\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_23\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_23\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_23\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_24\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_24\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_24\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_24\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_24\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_24\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_24\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_24\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_24\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_24\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_24\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_24\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_24\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_24\:Poor_Quality = "2" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_24\:Poor_Quality_Retrieved = "2" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_24\:Poor_Quality_Retrieved_Average_Sigma = "2.113266" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_25\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_25\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_25\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_25\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_25\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_25\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_25\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_25\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_25\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_25\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_25\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_25\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_25\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_25\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_25\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_25\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_26\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_26\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_26\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_26\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_26\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_26\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_26\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_26\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_26\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_26\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_26\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_26\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_26\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_26\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_26\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:LOQC\:Quality_Record_26\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:SIQ\:Grid_Point_Type = "Sea_Ice" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:SIQ\:SSS_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:SIQ\:SST_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:SIQ\:WS_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:SIQ\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:SIQ\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:SIQ\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:SIQ\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:SIQ\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:SIQ\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:SIQ\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:SIQ\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:SIQ\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:SIQ\:Poor_Quality = "64" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:SIQ\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_0\:SIQ\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:Retrieval_Scheme = "2" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:Land_Rejected = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:Too_Close_To_Land_Rejected = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:Ice_Rejected = "10855" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:Missing_ECMWF_Rejected = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:Too_Few_Measurements_Rejected = "18084" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:Good_Quality_Grid_Points = "29636" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:Poor_Quality_Grid_Points = "4896" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:SQ\:Grid_Point_Type = "Sea" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:SQ\:SSS_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:SQ\:SST_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:SQ\:WS_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:SQ\:Good_Quality = "23293" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:SQ\:Good_Quality_Retrieved = "16753" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:SQ\:Good_Quality_Retrieved_Average_Sigma = "2.016282" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:SQ\:Good_Quality_Failed_Outside_Valid_Range = "78" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:SQ\:Good_Quality_Failed_Sigma_Too_High = "479" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:SQ\:Good_Quality_Failed_Poor_Fit = "5999" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:SQ\:Good_Quality_Failed_Marquardt = "4" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:SQ\:Good_Quality_Failed_Maxiter = "273" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:SQ\:Good_Quality_Failed_OOLUT = "555" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:SQ\:Poor_Quality = "2426" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:SQ\:Poor_Quality_Retrieved = "1638" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:SQ\:Poor_Quality_Retrieved_Average_Sigma = "2.984403" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:NCQ\:Grid_Point_Type = "Near_Coast" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:NCQ\:SSS_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:NCQ\:SST_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:NCQ\:WS_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:NCQ\:Good_Quality = "6343" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:NCQ\:Good_Quality_Retrieved = "2879" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:NCQ\:Good_Quality_Retrieved_Average_Sigma = "1.380678" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:NCQ\:Good_Quality_Failed_Outside_Valid_Range = "281" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:NCQ\:Good_Quality_Failed_Sigma_Too_High = "532" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:NCQ\:Good_Quality_Failed_Poor_Fit = "3163" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:NCQ\:Good_Quality_Failed_Marquardt = "167" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:NCQ\:Good_Quality_Failed_Maxiter = "402" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:NCQ\:Good_Quality_Failed_OOLUT = "818" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:NCQ\:Poor_Quality = "2470" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:NCQ\:Poor_Quality_Retrieved = "1286" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:NCQ\:Poor_Quality_Retrieved_Average_Sigma = "1.503417" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_0\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_0\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_0\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_0\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_0\:Good_Quality = "559" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_0\:Good_Quality_Retrieved = "130" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_0\:Good_Quality_Retrieved_Average_Sigma = "1.956271" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_0\:Good_Quality_Failed_Outside_Valid_Range = "189" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_0\:Good_Quality_Failed_Sigma_Too_High = "265" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_0\:Good_Quality_Failed_Poor_Fit = "323" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_0\:Good_Quality_Failed_Marquardt = "121" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_0\:Good_Quality_Failed_Maxiter = "121" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_0\:Good_Quality_Failed_OOLUT = "326" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_0\:Poor_Quality = "106" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_0\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_0\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_1\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_1\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_1\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_1\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_1\:Good_Quality = "486" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_1\:Good_Quality_Retrieved = "228" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_1\:Good_Quality_Retrieved_Average_Sigma = "2.158294" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_1\:Good_Quality_Failed_Outside_Valid_Range = "59" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_1\:Good_Quality_Failed_Sigma_Too_High = "85" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_1\:Good_Quality_Failed_Poor_Fit = "245" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_1\:Good_Quality_Failed_Marquardt = "36" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_1\:Good_Quality_Failed_Maxiter = "40" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_1\:Good_Quality_Failed_OOLUT = "136" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_1\:Poor_Quality = "233" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_1\:Poor_Quality_Retrieved = "13" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_1\:Poor_Quality_Retrieved_Average_Sigma = "4.621669" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_2\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_2\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_2\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_2\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_2\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_2\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_2\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_2\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_2\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_2\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_2\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_2\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_2\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_2\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_2\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_2\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_3\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_3\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_3\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_3\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_3\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_3\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_3\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_3\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_3\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_3\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_3\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_3\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_3\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_3\:Poor_Quality = "3" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_3\:Poor_Quality_Retrieved = "1" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_3\:Poor_Quality_Retrieved_Average_Sigma = "2.825164" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_4\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_4\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_4\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_4\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_4\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_4\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_4\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_4\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_4\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_4\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_4\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_4\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_4\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_4\:Poor_Quality = "233" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_4\:Poor_Quality_Retrieved = "182" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_4\:Poor_Quality_Retrieved_Average_Sigma = "4.031709" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_5\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_5\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_5\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_5\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_5\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_5\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_5\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_5\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_5\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_5\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_5\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_5\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_5\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_5\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_5\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_5\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_6\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_6\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_6\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_6\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_6\:Good_Quality = "16" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_6\:Good_Quality_Retrieved = "14" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_6\:Good_Quality_Retrieved_Average_Sigma = "1.316742" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_6\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_6\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_6\:Good_Quality_Failed_Poor_Fit = "2" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_6\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_6\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_6\:Good_Quality_Failed_OOLUT = "1" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_6\:Poor_Quality = "22" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_6\:Poor_Quality_Retrieved = "16" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_6\:Poor_Quality_Retrieved_Average_Sigma = "1.820999" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_7\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_7\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_7\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_7\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_7\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_7\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_7\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_7\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_7\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_7\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_7\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_7\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_7\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_7\:Poor_Quality = "113" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_7\:Poor_Quality_Retrieved = "48" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_7\:Poor_Quality_Retrieved_Average_Sigma = "1.882463" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_8\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_8\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_8\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_8\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_8\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_8\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_8\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_8\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_8\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_8\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_8\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_8\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_8\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_8\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_8\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_8\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_9\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_9\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_9\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_9\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_9\:Good_Quality = "1485" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_9\:Good_Quality_Retrieved = "821" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_9\:Good_Quality_Retrieved_Average_Sigma = "2.183326" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_9\:Good_Quality_Failed_Outside_Valid_Range = "2" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_9\:Good_Quality_Failed_Sigma_Too_High = "57" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_9\:Good_Quality_Failed_Poor_Fit = "544" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_9\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_9\:Good_Quality_Failed_Maxiter = "247" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_9\:Good_Quality_Failed_OOLUT = "194" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_9\:Poor_Quality = "11" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_9\:Poor_Quality_Retrieved = "1" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_9\:Poor_Quality_Retrieved_Average_Sigma = "4.586421" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_10\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_10\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_10\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_10\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_10\:Good_Quality = "6940" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_10\:Good_Quality_Retrieved = "4685" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_10\:Good_Quality_Retrieved_Average_Sigma = "2.610784" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_10\:Good_Quality_Failed_Outside_Valid_Range = "102" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_10\:Good_Quality_Failed_Sigma_Too_High = "601" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_10\:Good_Quality_Failed_Poor_Fit = "1779" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_10\:Good_Quality_Failed_Marquardt = "14" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_10\:Good_Quality_Failed_Maxiter = "71" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_10\:Good_Quality_Failed_OOLUT = "604" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_10\:Poor_Quality = "508" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_10\:Poor_Quality_Retrieved = "216" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_10\:Poor_Quality_Retrieved_Average_Sigma = "4.321773" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_11\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_11\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_11\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_11\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_11\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_11\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_11\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_11\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_11\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_11\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_11\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_11\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_11\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_11\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_11\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_11\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_12\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_12\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_12\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_12\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_12\:Good_Quality = "232" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_12\:Good_Quality_Retrieved = "154" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_12\:Good_Quality_Retrieved_Average_Sigma = "1.546095" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_12\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_12\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_12\:Good_Quality_Failed_Poor_Fit = "73" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_12\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_12\:Good_Quality_Failed_Maxiter = "5" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_12\:Good_Quality_Failed_OOLUT = "17" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_12\:Poor_Quality = "55" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_12\:Poor_Quality_Retrieved = "44" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_12\:Poor_Quality_Retrieved_Average_Sigma = "2.515923" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_13\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_13\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_13\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_13\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_13\:Good_Quality = "11990" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_13\:Good_Quality_Retrieved = "9022" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_13\:Good_Quality_Retrieved_Average_Sigma = "2.096603" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_13\:Good_Quality_Failed_Outside_Valid_Range = "7" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_13\:Good_Quality_Failed_Sigma_Too_High = "3" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_13\:Good_Quality_Failed_Poor_Fit = "2966" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_13\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_13\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_13\:Good_Quality_Failed_OOLUT = "58" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_13\:Poor_Quality = "997" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_13\:Poor_Quality_Retrieved = "849" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_13\:Poor_Quality_Retrieved_Average_Sigma = "3.150212" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_14\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_14\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_14\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_14\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_14\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_14\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_14\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_14\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_14\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_14\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_14\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_14\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_14\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_14\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_14\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_14\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_15\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_15\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_15\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_15\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_15\:Good_Quality = "830" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_15\:Good_Quality_Retrieved = "539" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_15\:Good_Quality_Retrieved_Average_Sigma = "1.062494" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_15\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_15\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_15\:Good_Quality_Failed_Poor_Fit = "288" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_15\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_15\:Good_Quality_Failed_Maxiter = "3" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_15\:Good_Quality_Failed_OOLUT = "13" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_15\:Poor_Quality = "1379" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_15\:Poor_Quality_Retrieved = "1021" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_15\:Poor_Quality_Retrieved_Average_Sigma = "1.095964" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_16\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_16\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_16\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_16\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_16\:Good_Quality = "7097" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_16\:Good_Quality_Retrieved = "4038" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_16\:Good_Quality_Retrieved_Average_Sigma = "0.801339" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_16\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_16\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_16\:Good_Quality_Failed_Poor_Fit = "2942" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_16\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_16\:Good_Quality_Failed_Maxiter = "188" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_16\:Good_Quality_Failed_OOLUT = "24" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_16\:Poor_Quality = "1043" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_16\:Poor_Quality_Retrieved = "438" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_16\:Poor_Quality_Retrieved_Average_Sigma = "1.589996" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_17\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_17\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_17\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_17\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_17\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_17\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_17\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_17\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_17\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_17\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_17\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_17\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_17\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_17\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_17\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_17\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_18\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_18\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_18\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_18\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_18\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_18\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_18\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_18\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_18\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_18\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_18\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_18\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_18\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_18\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_18\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_18\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_19\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_19\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_19\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_19\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_19\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_19\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_19\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_19\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_19\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_19\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_19\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_19\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_19\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_19\:Poor_Quality = "141" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_19\:Poor_Quality_Retrieved = "52" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_19\:Poor_Quality_Retrieved_Average_Sigma = "4.370056" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_20\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_20\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_20\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_20\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_20\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_20\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_20\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_20\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_20\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_20\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_20\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_20\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_20\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_20\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_20\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_20\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_21\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_21\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_21\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_21\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_21\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_21\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_21\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_21\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_21\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_21\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_21\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_21\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_21\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_21\:Poor_Quality = "8" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_21\:Poor_Quality_Retrieved = "5" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_21\:Poor_Quality_Retrieved_Average_Sigma = "2.781770" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_22\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_22\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_22\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_22\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_22\:Good_Quality = "1" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_22\:Good_Quality_Retrieved = "1" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_22\:Good_Quality_Retrieved_Average_Sigma = "2.728715" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_22\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_22\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_22\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_22\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_22\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_22\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_22\:Poor_Quality = "42" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_22\:Poor_Quality_Retrieved = "36" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_22\:Poor_Quality_Retrieved_Average_Sigma = "3.373684" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_23\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_23\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_23\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_23\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_23\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_23\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_23\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_23\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_23\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_23\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_23\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_23\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_23\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_23\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_23\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_23\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_24\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_24\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_24\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_24\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_24\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_24\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_24\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_24\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_24\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_24\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_24\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_24\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_24\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_24\:Poor_Quality = "2" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_24\:Poor_Quality_Retrieved = "2" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_24\:Poor_Quality_Retrieved_Average_Sigma = "2.176347" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_25\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_25\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_25\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_25\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_25\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_25\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_25\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_25\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_25\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_25\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_25\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_25\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_25\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_25\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_25\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_25\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_26\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_26\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_26\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_26\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_26\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_26\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_26\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_26\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_26\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_26\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_26\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_26\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_26\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_26\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_26\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:LOQC\:Quality_Record_26\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:SIQ\:Grid_Point_Type = "Sea_Ice" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:SIQ\:SSS_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:SIQ\:SST_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:SIQ\:WS_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:SIQ\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:SIQ\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:SIQ\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:SIQ\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:SIQ\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:SIQ\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:SIQ\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:SIQ\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:SIQ\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:SIQ\:Poor_Quality = "64" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:SIQ\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_1\:SIQ\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:Retrieval_Scheme = "3" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:Land_Rejected = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:Too_Close_To_Land_Rejected = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:Ice_Rejected = "10855" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:Missing_ECMWF_Rejected = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:Too_Few_Measurements_Rejected = "18084" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:Good_Quality_Grid_Points = "29636" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:Poor_Quality_Grid_Points = "4896" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:SQ\:Grid_Point_Type = "Sea" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:SQ\:SSS_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:SQ\:SST_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:SQ\:WS_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:SQ\:Good_Quality = "23293" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:SQ\:Good_Quality_Retrieved = "17816" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:SQ\:Good_Quality_Retrieved_Average_Sigma = "1.959542" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:SQ\:Good_Quality_Failed_Outside_Valid_Range = "81" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:SQ\:Good_Quality_Failed_Sigma_Too_High = "478" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:SQ\:Good_Quality_Failed_Poor_Fit = "5037" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:SQ\:Good_Quality_Failed_Marquardt = "4" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:SQ\:Good_Quality_Failed_Maxiter = "110" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:SQ\:Good_Quality_Failed_OOLUT = "555" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:SQ\:Poor_Quality = "2426" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:SQ\:Poor_Quality_Retrieved = "1661" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:SQ\:Poor_Quality_Retrieved_Average_Sigma = "2.933723" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:NCQ\:Grid_Point_Type = "Near_Coast" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:NCQ\:SSS_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:NCQ\:SST_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:NCQ\:WS_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:NCQ\:Good_Quality = "6343" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:NCQ\:Good_Quality_Retrieved = "3803" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:NCQ\:Good_Quality_Retrieved_Average_Sigma = "1.253443" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:NCQ\:Good_Quality_Failed_Outside_Valid_Range = "276" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:NCQ\:Good_Quality_Failed_Sigma_Too_High = "522" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:NCQ\:Good_Quality_Failed_Poor_Fit = "2247" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:NCQ\:Good_Quality_Failed_Marquardt = "152" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:NCQ\:Good_Quality_Failed_Maxiter = "411" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:NCQ\:Good_Quality_Failed_OOLUT = "773" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:NCQ\:Poor_Quality = "2470" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:NCQ\:Poor_Quality_Retrieved = "1367" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:NCQ\:Poor_Quality_Retrieved_Average_Sigma = "1.480500" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_0\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_0\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_0\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_0\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_0\:Good_Quality = "559" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_0\:Good_Quality_Retrieved = "131" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_0\:Good_Quality_Retrieved_Average_Sigma = "1.985529" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_0\:Good_Quality_Failed_Outside_Valid_Range = "183" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_0\:Good_Quality_Failed_Sigma_Too_High = "261" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_0\:Good_Quality_Failed_Poor_Fit = "325" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_0\:Good_Quality_Failed_Marquardt = "112" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_0\:Good_Quality_Failed_Maxiter = "130" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_0\:Good_Quality_Failed_OOLUT = "326" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_0\:Poor_Quality = "106" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_0\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_0\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_1\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_1\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_1\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_1\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_1\:Good_Quality = "486" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_1\:Good_Quality_Retrieved = "229" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_1\:Good_Quality_Retrieved_Average_Sigma = "2.167454" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_1\:Good_Quality_Failed_Outside_Valid_Range = "60" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_1\:Good_Quality_Failed_Sigma_Too_High = "82" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_1\:Good_Quality_Failed_Poor_Fit = "244" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_1\:Good_Quality_Failed_Marquardt = "30" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_1\:Good_Quality_Failed_Maxiter = "45" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_1\:Good_Quality_Failed_OOLUT = "135" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_1\:Poor_Quality = "233" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_1\:Poor_Quality_Retrieved = "13" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_1\:Poor_Quality_Retrieved_Average_Sigma = "4.597799" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_2\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_2\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_2\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_2\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_2\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_2\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_2\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_2\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_2\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_2\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_2\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_2\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_2\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_2\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_2\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_2\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_3\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_3\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_3\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_3\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_3\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_3\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_3\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_3\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_3\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_3\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_3\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_3\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_3\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_3\:Poor_Quality = "3" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_3\:Poor_Quality_Retrieved = "1" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_3\:Poor_Quality_Retrieved_Average_Sigma = "2.726585" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_4\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_4\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_4\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_4\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_4\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_4\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_4\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_4\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_4\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_4\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_4\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_4\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_4\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_4\:Poor_Quality = "233" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_4\:Poor_Quality_Retrieved = "182" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_4\:Poor_Quality_Retrieved_Average_Sigma = "3.945308" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_5\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_5\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_5\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_5\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_5\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_5\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_5\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_5\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_5\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_5\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_5\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_5\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_5\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_5\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_5\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_5\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_6\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_6\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_6\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_6\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_6\:Good_Quality = "16" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_6\:Good_Quality_Retrieved = "14" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_6\:Good_Quality_Retrieved_Average_Sigma = "1.307737" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_6\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_6\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_6\:Good_Quality_Failed_Poor_Fit = "2" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_6\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_6\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_6\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_6\:Poor_Quality = "22" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_6\:Poor_Quality_Retrieved = "19" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_6\:Poor_Quality_Retrieved_Average_Sigma = "1.902701" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_7\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_7\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_7\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_7\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_7\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_7\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_7\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_7\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_7\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_7\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_7\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_7\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_7\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_7\:Poor_Quality = "113" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_7\:Poor_Quality_Retrieved = "58" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_7\:Poor_Quality_Retrieved_Average_Sigma = "1.925949" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_8\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_8\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_8\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_8\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_8\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_8\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_8\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_8\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_8\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_8\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_8\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_8\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_8\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_8\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_8\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_8\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_9\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_9\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_9\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_9\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_9\:Good_Quality = "1485" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_9\:Good_Quality_Retrieved = "825" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_9\:Good_Quality_Retrieved_Average_Sigma = "2.191673" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_9\:Good_Quality_Failed_Outside_Valid_Range = "1" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_9\:Good_Quality_Failed_Sigma_Too_High = "54" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_9\:Good_Quality_Failed_Poor_Fit = "544" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_9\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_9\:Good_Quality_Failed_Maxiter = "247" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_9\:Good_Quality_Failed_OOLUT = "190" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_9\:Poor_Quality = "11" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_9\:Poor_Quality_Retrieved = "1" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_9\:Poor_Quality_Retrieved_Average_Sigma = "4.534814" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_10\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_10\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_10\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_10\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_10\:Good_Quality = "6940" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_10\:Good_Quality_Retrieved = "4685" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_10\:Good_Quality_Retrieved_Average_Sigma = "2.611991" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_10\:Good_Quality_Failed_Outside_Valid_Range = "102" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_10\:Good_Quality_Failed_Sigma_Too_High = "600" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_10\:Good_Quality_Failed_Poor_Fit = "1779" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_10\:Good_Quality_Failed_Marquardt = "14" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_10\:Good_Quality_Failed_Maxiter = "72" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_10\:Good_Quality_Failed_OOLUT = "603" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_10\:Poor_Quality = "508" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_10\:Poor_Quality_Retrieved = "218" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_10\:Poor_Quality_Retrieved_Average_Sigma = "4.334874" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_11\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_11\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_11\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_11\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_11\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_11\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_11\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_11\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_11\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_11\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_11\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_11\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_11\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_11\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_11\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_11\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_12\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_12\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_12\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_12\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_12\:Good_Quality = "232" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_12\:Good_Quality_Retrieved = "156" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_12\:Good_Quality_Retrieved_Average_Sigma = "1.521774" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_12\:Good_Quality_Failed_Outside_Valid_Range = "1" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_12\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_12\:Good_Quality_Failed_Poor_Fit = "70" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_12\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_12\:Good_Quality_Failed_Maxiter = "7" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_12\:Good_Quality_Failed_OOLUT = "17" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_12\:Poor_Quality = "55" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_12\:Poor_Quality_Retrieved = "42" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_12\:Poor_Quality_Retrieved_Average_Sigma = "2.482193" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_13\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_13\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_13\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_13\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_13\:Good_Quality = "11990" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_13\:Good_Quality_Retrieved = "9532" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_13\:Good_Quality_Retrieved_Average_Sigma = "2.064730" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_13\:Good_Quality_Failed_Outside_Valid_Range = "10" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_13\:Good_Quality_Failed_Sigma_Too_High = "3" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_13\:Good_Quality_Failed_Poor_Fit = "2454" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_13\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_13\:Good_Quality_Failed_Maxiter = "1" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_13\:Good_Quality_Failed_OOLUT = "42" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_13\:Poor_Quality = "997" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_13\:Poor_Quality_Retrieved = "857" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_13\:Poor_Quality_Retrieved_Average_Sigma = "3.092174" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_14\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_14\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_14\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_14\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_14\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_14\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_14\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_14\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_14\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_14\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_14\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_14\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_14\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_14\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_14\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_14\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_15\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_15\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_15\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_15\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_15\:Good_Quality = "830" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_15\:Good_Quality_Retrieved = "677" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_15\:Good_Quality_Retrieved_Average_Sigma = "1.047869" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_15\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_15\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_15\:Good_Quality_Failed_Poor_Fit = "153" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_15\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_15\:Good_Quality_Failed_Maxiter = "1" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_15\:Good_Quality_Failed_OOLUT = "4" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_15\:Poor_Quality = "1379" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_15\:Poor_Quality_Retrieved = "1092" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_15\:Poor_Quality_Retrieved_Average_Sigma = "1.087475" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_16\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_16\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_16\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_16\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_16\:Good_Quality = "7097" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_16\:Good_Quality_Retrieved = "5369" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_16\:Good_Quality_Retrieved_Average_Sigma = "0.787403" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_16\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_16\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_16\:Good_Quality_Failed_Poor_Fit = "1713" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_16\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_16\:Good_Quality_Failed_Maxiter = "18" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_16\:Good_Quality_Failed_OOLUT = "11" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_16\:Poor_Quality = "1043" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_16\:Poor_Quality_Retrieved = "450" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_16\:Poor_Quality_Retrieved_Average_Sigma = "1.581808" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_17\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_17\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_17\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_17\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_17\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_17\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_17\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_17\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_17\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_17\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_17\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_17\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_17\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_17\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_17\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_17\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_18\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_18\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_18\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_18\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_18\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_18\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_18\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_18\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_18\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_18\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_18\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_18\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_18\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_18\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_18\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_18\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_19\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_19\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_19\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_19\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_19\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_19\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_19\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_19\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_19\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_19\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_19\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_19\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_19\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_19\:Poor_Quality = "141" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_19\:Poor_Quality_Retrieved = "51" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_19\:Poor_Quality_Retrieved_Average_Sigma = "4.372903" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_20\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_20\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_20\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_20\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_20\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_20\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_20\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_20\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_20\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_20\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_20\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_20\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_20\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_20\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_20\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_20\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_21\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_21\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_21\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_21\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_21\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_21\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_21\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_21\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_21\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_21\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_21\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_21\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_21\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_21\:Poor_Quality = "8" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_21\:Poor_Quality_Retrieved = "5" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_21\:Poor_Quality_Retrieved_Average_Sigma = "2.769263" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_22\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_22\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_22\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_22\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_22\:Good_Quality = "1" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_22\:Good_Quality_Retrieved = "1" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_22\:Good_Quality_Retrieved_Average_Sigma = "2.597888" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_22\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_22\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_22\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_22\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_22\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_22\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_22\:Poor_Quality = "42" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_22\:Poor_Quality_Retrieved = "37" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_22\:Poor_Quality_Retrieved_Average_Sigma = "3.355307" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_23\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_23\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_23\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_23\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_23\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_23\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_23\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_23\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_23\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_23\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_23\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_23\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_23\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_23\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_23\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_23\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_24\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_24\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_24\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_24\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_24\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_24\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_24\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_24\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_24\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_24\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_24\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_24\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_24\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_24\:Poor_Quality = "2" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_24\:Poor_Quality_Retrieved = "2" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_24\:Poor_Quality_Retrieved_Average_Sigma = "2.113266" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_25\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_25\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_25\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_25\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_25\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_25\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_25\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_25\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_25\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_25\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_25\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_25\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_25\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_25\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_25\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_25\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_26\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_26\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_26\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_26\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_26\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_26\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_26\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_26\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_26\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_26\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_26\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_26\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_26\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_26\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_26\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:LOQC\:Quality_Record_26\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:SIQ\:Grid_Point_Type = "Sea_Ice" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:SIQ\:SSS_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:SIQ\:SST_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:SIQ\:WS_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:SIQ\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:SIQ\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:SIQ\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:SIQ\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:SIQ\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:SIQ\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:SIQ\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:SIQ\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:SIQ\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:SIQ\:Poor_Quality = "64" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:SIQ\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_2\:SIQ\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:Retrieval_Scheme = "4" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:Land_Rejected = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:Too_Close_To_Land_Rejected = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:Ice_Rejected = "10855" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:Missing_ECMWF_Rejected = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:Too_Few_Measurements_Rejected = "18084" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:Good_Quality_Grid_Points = "29899" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:Poor_Quality_Grid_Points = "4633" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:SQ\:Grid_Point_Type = "Sea" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:SQ\:SSS_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:SQ\:SST_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:SQ\:WS_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:SQ\:Good_Quality = "23293" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:SQ\:Good_Quality_Retrieved = "21547" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:SQ\:Good_Quality_Retrieved_Average_Sigma = "0.736739" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:SQ\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:SQ\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:SQ\:Good_Quality_Failed_Poor_Fit = "1746" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:SQ\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:SQ\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:SQ\:Good_Quality_Failed_OOLUT = "1638" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:SQ\:Poor_Quality = "2426" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:SQ\:Poor_Quality_Retrieved = "1988" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:SQ\:Poor_Quality_Retrieved_Average_Sigma = "1.498341" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:NCQ\:Grid_Point_Type = "Near_Coast" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:NCQ\:SSS_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:NCQ\:SST_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:NCQ\:WS_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:NCQ\:Good_Quality = "6606" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:NCQ\:Good_Quality_Retrieved = "5264" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:NCQ\:Good_Quality_Retrieved_Average_Sigma = "0.828990" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:NCQ\:Good_Quality_Failed_Outside_Valid_Range = "254" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:NCQ\:Good_Quality_Failed_Sigma_Too_High = "32" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:NCQ\:Good_Quality_Failed_Poor_Fit = "1330" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:NCQ\:Good_Quality_Failed_Marquardt = "8" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:NCQ\:Good_Quality_Failed_Maxiter = "2" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:NCQ\:Good_Quality_Failed_OOLUT = "927" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:NCQ\:Poor_Quality = "2207" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:NCQ\:Poor_Quality_Retrieved = "1429" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:NCQ\:Poor_Quality_Retrieved_Average_Sigma = "1.448753" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_0\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_0\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_0\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_0\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_0\:Good_Quality = "559" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_0\:Good_Quality_Retrieved = "358" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_0\:Good_Quality_Retrieved_Average_Sigma = "0.674638" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_0\:Good_Quality_Failed_Outside_Valid_Range = "30" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_0\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_0\:Good_Quality_Failed_Poor_Fit = "190" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_0\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_0\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_0\:Good_Quality_Failed_OOLUT = "201" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_0\:Poor_Quality = "106" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_0\:Poor_Quality_Retrieved = "29" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_0\:Poor_Quality_Retrieved_Average_Sigma = "1.338563" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_1\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_1\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_1\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_1\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_1\:Good_Quality = "486" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_1\:Good_Quality_Retrieved = "385" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_1\:Good_Quality_Retrieved_Average_Sigma = "0.616946" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_1\:Good_Quality_Failed_Outside_Valid_Range = "4" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_1\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_1\:Good_Quality_Failed_Poor_Fit = "101" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_1\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_1\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_1\:Good_Quality_Failed_OOLUT = "101" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_1\:Poor_Quality = "233" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_1\:Poor_Quality_Retrieved = "136" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_1\:Poor_Quality_Retrieved_Average_Sigma = "1.539670" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_2\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_2\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_2\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_2\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_2\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_2\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_2\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_2\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_2\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_2\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_2\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_2\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_2\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_2\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_2\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_2\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_3\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_3\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_3\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_3\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_3\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_3\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_3\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_3\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_3\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_3\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_3\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_3\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_3\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_3\:Poor_Quality = "3" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_3\:Poor_Quality_Retrieved = "1" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_3\:Poor_Quality_Retrieved_Average_Sigma = "2.143224" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_4\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_4\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_4\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_4\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_4\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_4\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_4\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_4\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_4\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_4\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_4\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_4\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_4\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_4\:Poor_Quality = "233" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_4\:Poor_Quality_Retrieved = "187" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_4\:Poor_Quality_Retrieved_Average_Sigma = "1.582498" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_5\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_5\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_5\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_5\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_5\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_5\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_5\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_5\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_5\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_5\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_5\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_5\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_5\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_5\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_5\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_5\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_6\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_6\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_6\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_6\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_6\:Good_Quality = "16" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_6\:Good_Quality_Retrieved = "15" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_6\:Good_Quality_Retrieved_Average_Sigma = "1.357438" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_6\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_6\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_6\:Good_Quality_Failed_Poor_Fit = "1" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_6\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_6\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_6\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_6\:Poor_Quality = "22" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_6\:Poor_Quality_Retrieved = "19" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_6\:Poor_Quality_Retrieved_Average_Sigma = "2.030221" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_7\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_7\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_7\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_7\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_7\:Good_Quality = "28" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_7\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_7\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_7\:Good_Quality_Failed_Outside_Valid_Range = "19" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_7\:Good_Quality_Failed_Sigma_Too_High = "4" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_7\:Good_Quality_Failed_Poor_Fit = "28" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_7\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_7\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_7\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_7\:Poor_Quality = "85" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_7\:Poor_Quality_Retrieved = "53" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_7\:Poor_Quality_Retrieved_Average_Sigma = "1.845069" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_8\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_8\:SSS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_8\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_8\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_8\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_8\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_8\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_8\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_8\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_8\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_8\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_8\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_8\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_8\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_8\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_8\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_9\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_9\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_9\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_9\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_9\:Good_Quality = "1485" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_9\:Good_Quality_Retrieved = "1275" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_9\:Good_Quality_Retrieved_Average_Sigma = "0.643317" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_9\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_9\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_9\:Good_Quality_Failed_Poor_Fit = "210" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_9\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_9\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_9\:Good_Quality_Failed_OOLUT = "210" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_9\:Poor_Quality = "11" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_9\:Poor_Quality_Retrieved = "6" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_9\:Poor_Quality_Retrieved_Average_Sigma = "1.393877" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_10\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_10\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_10\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_10\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_10\:Good_Quality = "6940" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_10\:Good_Quality_Retrieved = "6223" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_10\:Good_Quality_Retrieved_Average_Sigma = "0.743647" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_10\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_10\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_10\:Good_Quality_Failed_Poor_Fit = "717" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_10\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_10\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_10\:Good_Quality_Failed_OOLUT = "717" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_10\:Poor_Quality = "508" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_10\:Poor_Quality_Retrieved = "387" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_10\:Poor_Quality_Retrieved_Average_Sigma = "1.451606" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_11\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_11\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_11\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_11\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_11\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_11\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_11\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_11\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_11\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_11\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_11\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_11\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_11\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_11\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_11\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_11\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_12\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_12\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_12\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_12\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_12\:Good_Quality = "232" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_12\:Good_Quality_Retrieved = "213" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_12\:Good_Quality_Retrieved_Average_Sigma = "0.741777" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_12\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_12\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_12\:Good_Quality_Failed_Poor_Fit = "19" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_12\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_12\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_12\:Good_Quality_Failed_OOLUT = "17" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_12\:Poor_Quality = "55" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_12\:Poor_Quality_Retrieved = "42" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_12\:Poor_Quality_Retrieved_Average_Sigma = "2.121626" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_13\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_13\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_13\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_13\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_13\:Good_Quality = "11990" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_13\:Good_Quality_Retrieved = "11136" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_13\:Good_Quality_Retrieved_Average_Sigma = "0.731001" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_13\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_13\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_13\:Good_Quality_Failed_Poor_Fit = "854" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_13\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_13\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_13\:Good_Quality_Failed_OOLUT = "813" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_13\:Poor_Quality = "997" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_13\:Poor_Quality_Retrieved = "847" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_13\:Poor_Quality_Retrieved_Average_Sigma = "1.560844" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_14\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_14\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_14\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_14\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_14\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_14\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_14\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_14\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_14\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_14\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_14\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_14\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_14\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_14\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_14\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_14\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_15\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_15\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_15\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_15\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_15\:Good_Quality = "830" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_15\:Good_Quality_Retrieved = "722" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_15\:Good_Quality_Retrieved_Average_Sigma = "1.117939" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_15\:Good_Quality_Failed_Outside_Valid_Range = "1" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_15\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_15\:Good_Quality_Failed_Poor_Fit = "107" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_15\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_15\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_15\:Good_Quality_Failed_OOLUT = "39" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_15\:Poor_Quality = "1379" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_15\:Poor_Quality_Retrieved = "1079" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_15\:Poor_Quality_Retrieved_Average_Sigma = "1.235114" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_16\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_16\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_16\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_16\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_16\:Good_Quality = "7332" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_16\:Good_Quality_Retrieved = "6483" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_16\:Good_Quality_Retrieved_Average_Sigma = "0.799682" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_16\:Good_Quality_Failed_Outside_Valid_Range = "200" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_16\:Good_Quality_Failed_Sigma_Too_High = "28" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_16\:Good_Quality_Failed_Poor_Fit = "849" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_16\:Good_Quality_Failed_Marquardt = "8" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_16\:Good_Quality_Failed_Maxiter = "2" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_16\:Good_Quality_Failed_OOLUT = "467" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_16\:Poor_Quality = "808" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_16\:Poor_Quality_Retrieved = "463" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_16\:Poor_Quality_Retrieved_Average_Sigma = "1.640629" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_17\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_17\:SSS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_17\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_17\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_17\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_17\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_17\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_17\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_17\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_17\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_17\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_17\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_17\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_17\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_17\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_17\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_18\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_18\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_18\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_18\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_18\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_18\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_18\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_18\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_18\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_18\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_18\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_18\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_18\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_18\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_18\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_18\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_19\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_19\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_19\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_19\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_19\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_19\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_19\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_19\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_19\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_19\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_19\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_19\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_19\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_19\:Poor_Quality = "141" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_19\:Poor_Quality_Retrieved = "127" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_19\:Poor_Quality_Retrieved_Average_Sigma = "1.663481" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_20\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_20\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_20\:SST_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_20\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_20\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_20\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_20\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_20\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_20\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_20\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_20\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_20\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_20\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_20\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_20\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_20\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_21\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_21\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_21\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_21\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_21\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_21\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_21\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_21\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_21\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_21\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_21\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_21\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_21\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_21\:Poor_Quality = "8" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_21\:Poor_Quality_Retrieved = "5" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_21\:Poor_Quality_Retrieved_Average_Sigma = "2.440643" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_22\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_22\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_22\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_22\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_22\:Good_Quality = "1" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_22\:Good_Quality_Retrieved = "1" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_22\:Good_Quality_Retrieved_Average_Sigma = "1.041794" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_22\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_22\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_22\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_22\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_22\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_22\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_22\:Poor_Quality = "42" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_22\:Poor_Quality_Retrieved = "36" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_22\:Poor_Quality_Retrieved_Average_Sigma = "1.924485" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_23\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_23\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_23\:SST_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_23\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_23\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_23\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_23\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_23\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_23\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_23\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_23\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_23\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_23\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_23\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_23\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_23\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_24\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_24\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_24\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_24\:WS_Class = "Low" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_24\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_24\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_24\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_24\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_24\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_24\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_24\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_24\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_24\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_24\:Poor_Quality = "2" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_24\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_24\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_25\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_25\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_25\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_25\:WS_Class = "Normal" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_25\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_25\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_25\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_25\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_25\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_25\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_25\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_25\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_25\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_25\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_25\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_25\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_26\:Grid_Point_Type = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_26\:SSS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_26\:SST_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_26\:WS_Class = "High" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_26\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_26\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_26\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_26\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_26\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_26\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_26\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_26\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_26\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_26\:Poor_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_26\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:LOQC\:Quality_Record_26\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:SIQ\:Grid_Point_Type = "Sea_Ice" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:SIQ\:SSS_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:SIQ\:SST_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:SIQ\:WS_Class = "All" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:SIQ\:Good_Quality = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:SIQ\:Good_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:SIQ\:Good_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:SIQ\:Good_Quality_Failed_Outside_Valid_Range = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:SIQ\:Good_Quality_Failed_Sigma_Too_High = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:SIQ\:Good_Quality_Failed_Poor_Fit = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:SIQ\:Good_Quality_Failed_Marquardt = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:SIQ\:Good_Quality_Failed_Maxiter = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:SIQ\:Good_Quality_Failed_OOLUT = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:SIQ\:Poor_Quality = "64" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:SIQ\:Poor_Quality_Retrieved = "0" ;
		string :VH\:SPH\:QI\:LORS\:Quality_Description_3\:SIQ\:Poor_Quality_Retrieved_Average_Sigma = "0.000000" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_0\:Retrieved_Parameter_0\:name = "SSS" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_0\:Retrieved_Parameter_0\:unit = "Practical Salinity Unit (PSU)" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_0\:Retrieved_Parameter_0\:description = "Surface salinity of the sea at gridpoint" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_0\:Retrieved_Parameter_1\:name = "SST" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_0\:Retrieved_Parameter_1\:unit = "Kelvin" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_0\:Retrieved_Parameter_1\:description = "Surface temperature of the sea at gridpoint" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_0\:Retrieved_Parameter_2\:name = "UN10" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_0\:Retrieved_Parameter_2\:unit = "m.s-1" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_0\:Retrieved_Parameter_2\:description = "U component of neutral wind 10m above surface" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_0\:Retrieved_Parameter_3\:name = "VN10" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_0\:Retrieved_Parameter_3\:unit = "m.s-1" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_0\:Retrieved_Parameter_3\:description = "V component of neutral wind 10m above surface" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_0\:Retrieved_Parameter_4\:name = "tec" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_0\:Retrieved_Parameter_4\:unit = "tecu" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_0\:Retrieved_Parameter_4\:description = "Total Electronic Content of the ionosphere below SMOS" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_0\:Retrieved_Parameter_5\:name = "not used" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_0\:Retrieved_Parameter_5\:unit = "none" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_0\:Retrieved_Parameter_5\:description = "no parameter defined" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_0\:Retrieved_Parameter_6\:name = "not used" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_0\:Retrieved_Parameter_6\:unit = "none" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_0\:Retrieved_Parameter_6\:description = "no parameter defined" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_0\:Retrieved_Parameter_7\:name = "not used" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_0\:Retrieved_Parameter_7\:unit = "none" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_0\:Retrieved_Parameter_7\:description = "no parameter defined" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_0\:Retrieved_Parameter_8\:name = "not used" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_0\:Retrieved_Parameter_8\:unit = "none" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_0\:Retrieved_Parameter_8\:description = "no parameter defined" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_0\:Retrieved_Parameter_9\:name = "not used" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_0\:Retrieved_Parameter_9\:unit = "none" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_0\:Retrieved_Parameter_9\:description = "no parameter defined" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_1\:Retrieved_Parameter_0\:name = "SSS" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_1\:Retrieved_Parameter_0\:unit = "Practical Salinity Unit (PSU)" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_1\:Retrieved_Parameter_0\:description = "Surface salinity of the sea at gridpoint" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_1\:Retrieved_Parameter_1\:name = "SST" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_1\:Retrieved_Parameter_1\:unit = "Kelvin" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_1\:Retrieved_Parameter_1\:description = "Surface temperature of the sea at gridpoint" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_1\:Retrieved_Parameter_2\:name = "UN10" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_1\:Retrieved_Parameter_2\:unit = "m.s-1" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_1\:Retrieved_Parameter_2\:description = "U component of neutral wind 10m above surface" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_1\:Retrieved_Parameter_3\:name = "VN10" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_1\:Retrieved_Parameter_3\:unit = "m.s-1" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_1\:Retrieved_Parameter_3\:description = "V component of neutral wind 10m above surface" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_1\:Retrieved_Parameter_4\:name = "tec" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_1\:Retrieved_Parameter_4\:unit = "tecu" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_1\:Retrieved_Parameter_4\:description = "Total Electronic Content of the ionosphere below SMOS" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_1\:Retrieved_Parameter_5\:name = "not used" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_1\:Retrieved_Parameter_5\:unit = "none" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_1\:Retrieved_Parameter_5\:description = "no parameter defined" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_1\:Retrieved_Parameter_6\:name = "not used" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_1\:Retrieved_Parameter_6\:unit = "none" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_1\:Retrieved_Parameter_6\:description = "no parameter defined" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_1\:Retrieved_Parameter_7\:name = "not used" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_1\:Retrieved_Parameter_7\:unit = "none" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_1\:Retrieved_Parameter_7\:description = "no parameter defined" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_1\:Retrieved_Parameter_8\:name = "not used" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_1\:Retrieved_Parameter_8\:unit = "none" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_1\:Retrieved_Parameter_8\:description = "no parameter defined" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_1\:Retrieved_Parameter_9\:name = "not used" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_1\:Retrieved_Parameter_9\:unit = "none" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_1\:Retrieved_Parameter_9\:description = "no parameter defined" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_2\:Retrieved_Parameter_0\:name = "SSS" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_2\:Retrieved_Parameter_0\:unit = "Practical Salinity Unit (PSU)" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_2\:Retrieved_Parameter_0\:description = "Surface salinity of the sea at gridpoint" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_2\:Retrieved_Parameter_1\:name = "SST" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_2\:Retrieved_Parameter_1\:unit = "Kelvin" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_2\:Retrieved_Parameter_1\:description = "Surface temperature of the sea at gridpoint" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_2\:Retrieved_Parameter_2\:name = "UN10" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_2\:Retrieved_Parameter_2\:unit = "m.s-1" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_2\:Retrieved_Parameter_2\:description = "U component of neutral wind 10m above surface" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_2\:Retrieved_Parameter_3\:name = "VN10" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_2\:Retrieved_Parameter_3\:unit = "m.s-1" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_2\:Retrieved_Parameter_3\:description = "V component of neutral wind 10m above surface" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_2\:Retrieved_Parameter_4\:name = "tec" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_2\:Retrieved_Parameter_4\:unit = "tecu" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_2\:Retrieved_Parameter_4\:description = "Total Electronic Content of the ionosphere below SMOS" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_2\:Retrieved_Parameter_5\:name = "not used" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_2\:Retrieved_Parameter_5\:unit = "none" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_2\:Retrieved_Parameter_5\:description = "no parameter defined" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_2\:Retrieved_Parameter_6\:name = "not used" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_2\:Retrieved_Parameter_6\:unit = "none" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_2\:Retrieved_Parameter_6\:description = "no parameter defined" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_2\:Retrieved_Parameter_7\:name = "not used" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_2\:Retrieved_Parameter_7\:unit = "none" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_2\:Retrieved_Parameter_7\:description = "no parameter defined" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_2\:Retrieved_Parameter_8\:name = "not used" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_2\:Retrieved_Parameter_8\:unit = "none" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_2\:Retrieved_Parameter_8\:description = "no parameter defined" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_2\:Retrieved_Parameter_9\:name = "not used" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_2\:Retrieved_Parameter_9\:unit = "none" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_2\:Retrieved_Parameter_9\:description = "no parameter defined" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_3\:Retrieved_Parameter_0\:name = "Acard" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_3\:Retrieved_Parameter_0\:unit = "dl" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_3\:Retrieved_Parameter_0\:description = "Acard coefficient for cardioid model" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_3\:Retrieved_Parameter_1\:name = "SST" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_3\:Retrieved_Parameter_1\:unit = "Kelvin" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_3\:Retrieved_Parameter_1\:description = "Surface temperature of the sea at gridpoint" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_3\:Retrieved_Parameter_2\:name = "not used" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_3\:Retrieved_Parameter_2\:unit = "none" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_3\:Retrieved_Parameter_2\:description = "no parameter defined" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_3\:Retrieved_Parameter_3\:name = "not used" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_3\:Retrieved_Parameter_3\:unit = "none" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_3\:Retrieved_Parameter_3\:description = "no parameter defined" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_3\:Retrieved_Parameter_4\:name = "not used" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_3\:Retrieved_Parameter_4\:unit = "none" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_3\:Retrieved_Parameter_4\:description = "no parameter defined" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_3\:Retrieved_Parameter_5\:name = "not used" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_3\:Retrieved_Parameter_5\:unit = "none" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_3\:Retrieved_Parameter_5\:description = "no parameter defined" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_3\:Retrieved_Parameter_6\:name = "not used" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_3\:Retrieved_Parameter_6\:unit = "none" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_3\:Retrieved_Parameter_6\:description = "no parameter defined" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_3\:Retrieved_Parameter_7\:name = "not used" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_3\:Retrieved_Parameter_7\:unit = "none" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_3\:Retrieved_Parameter_7\:description = "no parameter defined" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_3\:Retrieved_Parameter_8\:name = "not used" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_3\:Retrieved_Parameter_8\:unit = "none" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_3\:Retrieved_Parameter_8\:description = "no parameter defined" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_3\:Retrieved_Parameter_9\:name = "not used" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_3\:Retrieved_Parameter_9\:unit = "none" ;
		string :VH\:SPH\:L2PD\:LOM\:List_of_Retrieved_Parameters_3\:Retrieved_Parameter_9\:description = "no parameter defined" ;
		string :VH\:SPH\:MI\:SPH_Descriptor = "MIR_OSUDP2_SPH" ;
		string :VH\:SPH\:MI\:Checksum = "0186172426" ;
		string :VH\:SPH\:MI\:Header_Schema = "HDR_SM_XXXX_MIR_OSUDP2_0400.xsd" ;
		string :VH\:SPH\:MI\:Datablock_Schema = "DBL_SM_XXXX_MIR_OSUDP2_0401.binXschema.xml" ;
		string :VH\:SPH\:MI\:Header_Size = "168617" ;
		string :VH\:SPH\:MI\:Datablock_Size = "00017615474" ;
		string :VH\:SPH\:MI\:HW_Identifier = "0002" ;
		string :VH\:SPH\:MI\:TI\:Precise_Validity_Start = "UTC=2021-06-30T21:59:10.071954" ;
		string :VH\:SPH\:MI\:TI\:Precise_Validity_Stop = "UTC=2021-06-30T22:52:30.511865" ;
		string :VH\:SPH\:MI\:TI\:Abs_Orbit_Start = "+61281" ;
		string :VH\:SPH\:MI\:TI\:Start_Time_ANX_T = "4283.930491" ;
		string :VH\:SPH\:MI\:TI\:Abs_Orbit_Stop = "+61282" ;
		string :VH\:SPH\:MI\:TI\:Stop_Time_ANX_T = "1479.892790" ;
		string :VH\:SPH\:MI\:TI\:UTC_at_ANX = "UTC=2021-06-30T20:47:46.141463" ;
		string :VH\:SPH\:MI\:TI\:Long_at_ANX = "+138.381497" ;
		string :VH\:SPH\:MI\:TI\:Ascending_Flag = "A" ;
		string :VH\:SPH\:MI\:TI\:Polarisation_Flag = "F" ;
		string :VH\:SPH\:LODS\:Data_Set_0\:DS_Name = "SSS_SWATH" ;
		string :VH\:SPH\:LODS\:Data_Set_0\:DS_Type = "M" ;
		string :VH\:SPH\:LODS\:Data_Set_0\:DS_Size = "0017615474" ;
		string :VH\:SPH\:LODS\:Data_Set_0\:DS_Offset = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_0\:Num_DSR = "0000092713" ;
		string :VH\:SPH\:LODS\:Data_Set_0\:DSR_Size = "00000190" ;
		string :VH\:SPH\:LODS\:Data_Set_0\:Byte_Order = "0123" ;
		string :VH\:SPH\:LODS\:Data_Set_1\:DS_Name = "L1C_OS_FILE" ;
		string :VH\:SPH\:LODS\:Data_Set_1\:DS_Type = "R" ;
		string :VH\:SPH\:LODS\:Data_Set_1\:DS_Size = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_1\:DS_Offset = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_1\:Ref_Filename = "SM_OPER_MIR_SCSF1C_20210630T215911_20210630T225230_724_001_1" ;
		string :VH\:SPH\:LODS\:Data_Set_1\:Num_DSR = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_1\:DSR_Size = "00000000" ;
		string :VH\:SPH\:LODS\:Data_Set_1\:Byte_Order = "0000" ;
		string :VH\:SPH\:LODS\:Data_Set_2\:DS_Name = "DGG_FILE" ;
		string :VH\:SPH\:LODS\:Data_Set_2\:DS_Type = "R" ;
		string :VH\:SPH\:LODS\:Data_Set_2\:DS_Size = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_2\:DS_Offset = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_2\:Ref_Filename = "SM_OPER_AUX_DGG____20050101T000000_20500101T000000_300_003_3" ;
		string :VH\:SPH\:LODS\:Data_Set_2\:Num_DSR = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_2\:DSR_Size = "00000000" ;
		string :VH\:SPH\:LODS\:Data_Set_2\:Byte_Order = "0000" ;
		string :VH\:SPH\:LODS\:Data_Set_3\:DS_Name = "IERS_BULLETIN_B_FILE" ;
		string :VH\:SPH\:LODS\:Data_Set_3\:DS_Type = "R" ;
		string :VH\:SPH\:LODS\:Data_Set_3\:DS_Size = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_3\:DS_Offset = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_3\:Ref_Filename = "SM_OPER_AUX_BULL_B_20210402T000000_20500101T000000_120_001_3" ;
		string :VH\:SPH\:LODS\:Data_Set_3\:Num_DSR = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_3\:DSR_Size = "00000000" ;
		string :VH\:SPH\:LODS\:Data_Set_3\:Byte_Order = "0000" ;
		string :VH\:SPH\:LODS\:Data_Set_4\:DS_Name = "BESTFITPLANE_FILE" ;
		string :VH\:SPH\:LODS\:Data_Set_4\:DS_Type = "R" ;
		string :VH\:SPH\:LODS\:Data_Set_4\:DS_Size = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_4\:DS_Offset = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_4\:Ref_Filename = "SM_OPER_AUX_BFP____20050101T000000_20500101T000000_340_004_3" ;
		string :VH\:SPH\:LODS\:Data_Set_4\:Num_DSR = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_4\:DSR_Size = "00000000" ;
		string :VH\:SPH\:LODS\:Data_Set_4\:Byte_Order = "0000" ;
		string :VH\:SPH\:LODS\:Data_Set_5\:DS_Name = "MISPOINTING_FILE" ;
		string :VH\:SPH\:LODS\:Data_Set_5\:DS_Type = "R" ;
		string :VH\:SPH\:LODS\:Data_Set_5\:DS_Size = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_5\:DS_Offset = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_5\:Ref_Filename = "SM_OPER_AUX_MISP___20050101T000000_20500101T000000_300_004_3" ;
		string :VH\:SPH\:LODS\:Data_Set_5\:Num_DSR = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_5\:DSR_Size = "00000000" ;
		string :VH\:SPH\:LODS\:Data_Set_5\:Byte_Order = "0000" ;
		string :VH\:SPH\:LODS\:Data_Set_6\:DS_Name = "ECMWF_FILE" ;
		string :VH\:SPH\:LODS\:Data_Set_6\:DS_Type = "R" ;
		string :VH\:SPH\:LODS\:Data_Set_6\:DS_Size = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_6\:DS_Offset = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_6\:Ref_Filename = "SM_OPER_AUX_ECMWF__20210630T215902_20210630T230542_318_001_3" ;
		string :VH\:SPH\:LODS\:Data_Set_6\:Num_DSR = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_6\:DSR_Size = "00000000" ;
		string :VH\:SPH\:LODS\:Data_Set_6\:Byte_Order = "0000" ;
		string :VH\:SPH\:LODS\:Data_Set_7\:DS_Name = "FLAT_SEA_FILE" ;
		string :VH\:SPH\:LODS\:Data_Set_7\:DS_Type = "R" ;
		string :VH\:SPH\:LODS\:Data_Set_7\:DS_Size = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_7\:DS_Offset = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_7\:Ref_Filename = "SM_OPER_AUX_FLTSEA_20050101T000000_20500101T000000_001_012_3" ;
		string :VH\:SPH\:LODS\:Data_Set_7\:Num_DSR = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_7\:DSR_Size = "00000000" ;
		string :VH\:SPH\:LODS\:Data_Set_7\:Byte_Order = "0000" ;
		string :VH\:SPH\:LODS\:Data_Set_8\:DS_Name = "ROUGHNESS_IPSL_FILE" ;
		string :VH\:SPH\:LODS\:Data_Set_8\:DS_Type = "R" ;
		string :VH\:SPH\:LODS\:Data_Set_8\:DS_Size = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_8\:DS_Offset = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_8\:Ref_Filename = "SM_OPER_AUX_RGHNS1_20050101T000000_20500101T000000_001_016_3" ;
		string :VH\:SPH\:LODS\:Data_Set_8\:Num_DSR = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_8\:DSR_Size = "00000000" ;
		string :VH\:SPH\:LODS\:Data_Set_8\:Byte_Order = "0000" ;
		string :VH\:SPH\:LODS\:Data_Set_9\:DS_Name = "ROUGHNESS_IFREMER_FILE" ;
		string :VH\:SPH\:LODS\:Data_Set_9\:DS_Type = "R" ;
		string :VH\:SPH\:LODS\:Data_Set_9\:DS_Size = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_9\:DS_Offset = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_9\:Ref_Filename = "SM_OPER_AUX_RGHNS2_20050101T000000_20500101T000000_001_013_3" ;
		string :VH\:SPH\:LODS\:Data_Set_9\:Num_DSR = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_9\:DSR_Size = "00000000" ;
		string :VH\:SPH\:LODS\:Data_Set_9\:Byte_Order = "0000" ;
		string :VH\:SPH\:LODS\:Data_Set_10\:DS_Name = "ROUGHNESS_ICM_CSIC_FILE" ;
		string :VH\:SPH\:LODS\:Data_Set_10\:DS_Type = "R" ;
		string :VH\:SPH\:LODS\:Data_Set_10\:DS_Size = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_10\:DS_Offset = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_10\:Ref_Filename = "SM_OPER_AUX_RGHNS3_20050101T000000_20500101T000000_001_016_3" ;
		string :VH\:SPH\:LODS\:Data_Set_10\:Num_DSR = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_10\:DSR_Size = "00000000" ;
		string :VH\:SPH\:LODS\:Data_Set_10\:Byte_Order = "0000" ;
		string :VH\:SPH\:LODS\:Data_Set_11\:DS_Name = "GALAXY_OS_FILE" ;
		string :VH\:SPH\:LODS\:Data_Set_11\:DS_Type = "R" ;
		string :VH\:SPH\:LODS\:Data_Set_11\:DS_Size = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_11\:DS_Offset = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_11\:Ref_Filename = "SM_OPER_AUX_GAL_OS_20050101T000000_20500101T000000_001_011_3" ;
		string :VH\:SPH\:LODS\:Data_Set_11\:Num_DSR = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_11\:DSR_Size = "00000000" ;
		string :VH\:SPH\:LODS\:Data_Set_11\:Byte_Order = "0000" ;
		string :VH\:SPH\:LODS\:Data_Set_12\:DS_Name = "GALAXY_2OS_FILE" ;
		string :VH\:SPH\:LODS\:Data_Set_12\:DS_Type = "R" ;
		string :VH\:SPH\:LODS\:Data_Set_12\:DS_Size = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_12\:DS_Offset = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_12\:Ref_Filename = "SM_OPER_AUX_GAL2OS_20050101T000000_20500101T000000_001_016_3" ;
		string :VH\:SPH\:LODS\:Data_Set_12\:Num_DSR = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_12\:DSR_Size = "00000000" ;
		string :VH\:SPH\:LODS\:Data_Set_12\:Byte_Order = "0000" ;
		string :VH\:SPH\:LODS\:Data_Set_13\:DS_Name = "SUNGLINT_FILE" ;
		string :VH\:SPH\:LODS\:Data_Set_13\:DS_Type = "R" ;
		string :VH\:SPH\:LODS\:Data_Set_13\:DS_Size = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_13\:DS_Offset = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_13\:Ref_Filename = "SM_OPER_AUX_SGLINT_20050101T000000_20500101T000000_001_012_3" ;
		string :VH\:SPH\:LODS\:Data_Set_13\:Num_DSR = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_13\:DSR_Size = "00000000" ;
		string :VH\:SPH\:LODS\:Data_Set_13\:Byte_Order = "0000" ;
		string :VH\:SPH\:LODS\:Data_Set_14\:DS_Name = "ATMOS_FILE" ;
		string :VH\:SPH\:LODS\:Data_Set_14\:DS_Type = "R" ;
		string :VH\:SPH\:LODS\:Data_Set_14\:DS_Size = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_14\:DS_Offset = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_14\:Ref_Filename = "SM_OPER_AUX_ATMOS__20050101T000000_20500101T000000_001_010_3" ;
		string :VH\:SPH\:LODS\:Data_Set_14\:Num_DSR = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_14\:DSR_Size = "00000000" ;
		string :VH\:SPH\:LODS\:Data_Set_14\:Byte_Order = "0000" ;
		string :VH\:SPH\:LODS\:Data_Set_15\:DS_Name = "DISTAN_FILE" ;
		string :VH\:SPH\:LODS\:Data_Set_15\:DS_Type = "R" ;
		string :VH\:SPH\:LODS\:Data_Set_15\:DS_Size = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_15\:DS_Offset = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_15\:Ref_Filename = "SM_OPER_AUX_DISTAN_20050101T000000_20500101T000000_001_011_3" ;
		string :VH\:SPH\:LODS\:Data_Set_15\:Num_DSR = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_15\:DSR_Size = "00000000" ;
		string :VH\:SPH\:LODS\:Data_Set_15\:Byte_Order = "0000" ;
		string :VH\:SPH\:LODS\:Data_Set_16\:DS_Name = "CLIMATOLOGY_SSS_FILE" ;
		string :VH\:SPH\:LODS\:Data_Set_16\:DS_Type = "R" ;
		string :VH\:SPH\:LODS\:Data_Set_16\:DS_Size = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_16\:DS_Offset = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_16\:Ref_Filename = "SM_OPER_AUX_SSS____20050101T000000_20500101T000000_001_014_3" ;
		string :VH\:SPH\:LODS\:Data_Set_16\:Num_DSR = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_16\:DSR_Size = "00000000" ;
		string :VH\:SPH\:LODS\:Data_Set_16\:Byte_Order = "0000" ;
		string :VH\:SPH\:LODS\:Data_Set_17\:DS_Name = "CLIMATOLOGY_SSSCLI_FILE" ;
		string :VH\:SPH\:LODS\:Data_Set_17\:DS_Type = "R" ;
		string :VH\:SPH\:LODS\:Data_Set_17\:DS_Size = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_17\:DS_Offset = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_17\:Ref_Filename = "SM_OPER_AUX_SSSCLI_20050101T000000_20500101T000000_001_002_3" ;
		string :VH\:SPH\:LODS\:Data_Set_17\:Num_DSR = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_17\:DSR_Size = "00000000" ;
		string :VH\:SPH\:LODS\:Data_Set_17\:Byte_Order = "0000" ;
		string :VH\:SPH\:LODS\:Data_Set_18\:DS_Name = "OCEAN_SALINITY_CONFIG_FILE" ;
		string :VH\:SPH\:LODS\:Data_Set_18\:DS_Type = "R" ;
		string :VH\:SPH\:LODS\:Data_Set_18\:DS_Size = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_18\:DS_Offset = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_18\:Ref_Filename = "SM_OPER_AUX_CNFOSF_20050101T000000_20500101T000000_001_032_3" ;
		string :VH\:SPH\:LODS\:Data_Set_18\:Num_DSR = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_18\:DSR_Size = "00000000" ;
		string :VH\:SPH\:LODS\:Data_Set_18\:Byte_Order = "0000" ;
		string :VH\:SPH\:LODS\:Data_Set_19\:DS_Name = "OTT1F_FILE" ;
		string :VH\:SPH\:LODS\:Data_Set_19\:DS_Type = "R" ;
		string :VH\:SPH\:LODS\:Data_Set_19\:DS_Size = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_19\:DS_Offset = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_19\:Ref_Filename = "SM_OPER_AUX_OTT1F__20210624T082406_20500101T000000_700_001_1" ;
		string :VH\:SPH\:LODS\:Data_Set_19\:Num_DSR = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_19\:DSR_Size = "00000000" ;
		string :VH\:SPH\:LODS\:Data_Set_19\:Byte_Order = "0000" ;
		string :VH\:SPH\:LODS\:Data_Set_20\:DS_Name = "OTT2F_FILE" ;
		string :VH\:SPH\:LODS\:Data_Set_20\:DS_Type = "R" ;
		string :VH\:SPH\:LODS\:Data_Set_20\:DS_Size = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_20\:DS_Offset = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_20\:Ref_Filename = "SM_OPER_AUX_OTT2F__20210624T082406_20500101T000000_700_001_1" ;
		string :VH\:SPH\:LODS\:Data_Set_20\:Num_DSR = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_20\:DSR_Size = "00000000" ;
		string :VH\:SPH\:LODS\:Data_Set_20\:Byte_Order = "0000" ;
		string :VH\:SPH\:LODS\:Data_Set_21\:DS_Name = "OTT3F_FILE" ;
		string :VH\:SPH\:LODS\:Data_Set_21\:DS_Type = "R" ;
		string :VH\:SPH\:LODS\:Data_Set_21\:DS_Size = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_21\:DS_Offset = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_21\:Ref_Filename = "SM_OPER_AUX_OTT3F__20210624T082406_20500101T000000_700_001_1" ;
		string :VH\:SPH\:LODS\:Data_Set_21\:Num_DSR = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_21\:DSR_Size = "00000000" ;
		string :VH\:SPH\:LODS\:Data_Set_21\:Byte_Order = "0000" ;
		string :VH\:SPH\:LODS\:Data_Set_22\:DS_Name = "DGGRFI_FILE" ;
		string :VH\:SPH\:LODS\:Data_Set_22\:DS_Type = "R" ;
		string :VH\:SPH\:LODS\:Data_Set_22\:DS_Size = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_22\:DS_Offset = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_22\:Ref_Filename = "SM_OPER_AUX_DGGRFI_20210629T000711_20500101T000000_600_001_1" ;
		string :VH\:SPH\:LODS\:Data_Set_22\:Num_DSR = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_22\:DSR_Size = "00000000" ;
		string :VH\:SPH\:LODS\:Data_Set_22\:Byte_Order = "0000" ;
		string :VH\:SPH\:LODS\:Data_Set_23\:DS_Name = "MIXED_SCENE_OTT_FILE" ;
		string :VH\:SPH\:LODS\:Data_Set_23\:DS_Type = "R" ;
		string :VH\:SPH\:LODS\:Data_Set_23\:DS_Size = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_23\:DS_Offset = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_23\:Ref_Filename = "SM_OPER_AUX_MSOTT__20050101T000000_20500101T000000_001_002_3" ;
		string :VH\:SPH\:LODS\:Data_Set_23\:Num_DSR = "0000000000" ;
		string :VH\:SPH\:LODS\:Data_Set_23\:DSR_Size = "00000000" ;
		string :VH\:SPH\:LODS\:Data_Set_23\:Byte_Order = "0000" ;
		string :VH\:SPH\:L2PL\:Start_Lat = "-075.538036" ;
		string :VH\:SPH\:L2PL\:Start_Long = "-094.410663" ;
		string :VH\:SPH\:L2PL\:Stop_Lat = "+081.601490" ;
		string :VH\:SPH\:L2PL\:Stop_Long = "+017.400949" ;
		string :VH\:SPH\:L2PL\:Mid_Lat = "-005.823823" ;
		string :VH\:SPH\:L2PL\:Mid_Lon = "+114.700199" ;
		string :VH\:SPH\:L2PL\:Southernmost_Latitude = "-063.270000" ;
		string :VH\:SPH\:L2PL\:Southernmost_Gridpoint_ID = "7240286" ;
		string :VH\:SPH\:L2PL\:Northernmost_Latitude = "+080.555000" ;
		string :VH\:SPH\:L2PL\:Northernmost_Gridpoint_ID = "4094657" ;
		string :VH\:SPH\:L2PL\:Easternmost_Longitude = "+148.524002" ;
		string :VH\:SPH\:L2PL\:Easternmost_Gridpoint_ID = "7243351" ;
		string :VH\:SPH\:L2PL\:Westernmost_Longitude = "+023.934000" ;
		string :VH\:SPH\:L2PL\:Westernmost_Gridpoint_ID = "4081389" ;
		string :VH\:MPH\:Ref_Doc = "SO-TN-IDR-GS-0006" ;
		string :VH\:MPH\:Acquisition_Station = "SVLD" ;
		string :VH\:MPH\:Processing_Centre = "ESAC" ;
		string :VH\:MPH\:Logical_Proc_Centre = "FPC" ;
		string :VH\:MPH\:Product_Confidence = "NOMINAL" ;
		string :VH\:MPH\:OI\:Phase = "+001" ;
		string :VH\:MPH\:OI\:Cycle = "+037" ;
		string :VH\:MPH\:OI\:Rel_Orbit = "+01161" ;
		string :VH\:MPH\:OI\:Abs_Orbit = "+61281" ;
		string :VH\:MPH\:OI\:OSV_TAI = "TAI=2021-06-30T21:58:37.000000" ;
		string :VH\:MPH\:OI\:OSV_UTC = "UTC=2021-06-30T21:58:00.000000" ;
		string :VH\:MPH\:OI\:OSV_UT1 = "UT1=2021-06-30T21:58:00.590000" ;
		string :VH\:MPH\:OI\:X_Position = "+0146839.075" ;
		string :VH\:MPH\:OI\:Y_Position = "-2215887.397" ;
		string :VH\:MPH\:OI\:Z_Position = "-6791787.132" ;
		string :VH\:MPH\:OI\:X_Velocity = "-4093.431900" ;
		string :VH\:MPH\:OI\:Y_Velocity = "+5989.437140" ;
		string :VH\:MPH\:OI\:Z_Velocity = "-2043.308610" ;
		string :VH\:MPH\:OI\:Vector_Source = "FP" ;
		:history = "Mon Oct  2 16:02:44 2023: ncks -d n_grid_points,100,92700,1800 -v SSS_corr,Sigma_SSS_corr,Latitude,Longitude,Mean_acq_time,Dg_quality_SSS_corr /scratch1/NCEPDEV/stmp4/Shastri.Paturi/forAndrew/gdas.20210701/00/SSS/SM_OPER_MIR_OSUDP2_20210630T215911_20210630T225230_700_001_1.nc sss_smos_2_sub.nc" ;
		:NCO = "netCDF Operators version 5.0.6 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco)" ;
data:

 Dg_quality_SSS_corr = _, _, _, _, _, _, _, _, 247, 300, _, _, 125, _, 131, 
    298, 92, 306, 116, _, 219, _, _, _, _, 57, 154, 210, _, _, _, 168, 128, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, 288, _, _, _, 472, _ ;

 Latitude = -76.151, -77.41, -74.643, -71.861, -64.609, -63.034, -64.906, 
    -63.205, -55.638, -54.537, -57.479, -58.616, -48.685, -51.452, -44.391, 
    -46.513, -40.182, -42.866, -35.332, -39.175, -37.132, -33.301, -28.93, 
    -25.44, -14.805, -13.467, -16.861, -14.725, -4.935, -4.42, -2.378, 
    -5.508, 2.697, -3.076, 1.48, 10.232, 11.234, 13.737, 16.148, 18.106, 
    22.444, 17.864, 51.638, 69.291, 74.944, 74.356, 77.42, 77.959, 71.973, 
    80.454, 76.93, 87.38 ;

 Longitude = -157.126, 177.916, -170.177, 165.449, 143.108, 138.427, 147.869, 
    148.091, 134.345, 123.998, 144.011, 120.997, 126.188, 137.108, 122.752, 
    131.805, 122.686, 131.029, 123.431, 131.595, 117.177, 115.688, 114.405, 
    114.364, 119.251, 116.545, 113.311, 122.324, 117.944, 115.496, 111.48, 
    110.942, 110.625, 108.663, 118.323, 113.515, 110.075, 108.134, 110.859, 
    107.175, 112.003, 116.105, 101.016, 82.105, 85.012, 60.59, 64.585, 
    51.372, 58.422, 86.772, 37.611, 56.383 ;

 Mean_acq_time = 7851.918, 7851.919, 7851.919, _, 7851.922, 7851.922, 
    7851.922, 7851.922, 7851.924, 7851.924, 7851.923, 7851.924, 7851.925, 
    7851.925, 7851.926, 7851.926, 7851.927, 7851.927, 7851.928, 7851.927, 
    7851.928, 7851.929, 7851.93, _, 7851.932, 7851.932, 7851.932, 7851.932, 
    7851.934, 7851.934, _, 7851.935, 7851.936, 7851.935, _, 7851.937, 
    7851.937, _, 7851.938, 7851.938, _, 7851.938, _, _, 7851.95, 7851.95, 
    7851.951, 7851.951, 7851.951, 7851.951, 7851.952, 7851.952 ;

 SSS_corr = _, _, _, _, _, _, _, _, 30.59692, 34.46416, _, _, 29.57378, 
    33.6181, 32.66331, 38.32122, 30.43209, 28.0537, 35.61701, _, 33.53222, _, 
    _, _, 32.95224, 33.26748, 34.88172, 34.5612, _, _, _, 32.28378, 31.75333, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, 31.5253, 31.22411, 0.9942121, _, 
    33.04895, _ ;

 Sigma_SSS_corr = _, _, _, _, _, _, _, _, 1.943289, 2.015971, _, _, 2.21241, 
    4.420088, 2.091019, 3.159312, 1.382608, 2.935465, 1.132476, _, 1.895663, 
    _, _, _, 0.6969603, 0.5503999, 0.8192711, 1.835188, _, _, _, 0.8325468, 
    0.6733742, _, _, _, _, _, _, _, _, _, _, _, _, _, 2.208032, 2.230621, 
    213.0026, _, 3.79549, _ ;
}
