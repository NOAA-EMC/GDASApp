netcdf prof.nc {
dimensions:
	Location = 218 ;
	nvars = 2 ;
variables:
	int Location(Location) ;
		Location:suggested_chunk_dim = 218LL ;
	float nvars(nvars) ;
		nvars:suggested_chunk_dim = 100LL ;

// global attributes:
		string :_ioda_layout = "ObsGroup" ;
		:_ioda_layout_version = 0 ;
		:nrecs = 20 ;
		:nvars = 2 ;
		:odb_version = 1LL ;
		:date_time = 2018041512 ;
		:nlocs = 218 ;
		:nobs = 436 ;
data:

 Location = 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
    0, 0, 0, 0 ;

 nvars = 0, 0 ;

group: MetaData {
  variables:
  	int64 dateTime(Location) ;
  		dateTime:_FillValue = -3732782400LL ;
  		string dateTime:units = "seconds since 2018-04-15T12:00:00Z" ;
  	string date_time(Location) ;
  		string date_time:_FillValue = "" ;
  	float depth(Location) ;
  		depth:_FillValue = 9.96921e+36f ;
  	float latitude(Location) ;
  		latitude:_FillValue = 9.96921e+36f ;
  	float longitude(Location) ;
  		longitude:_FillValue = 9.96921e+36f ;
  	int sequenceNumber(Location) ;
  		sequenceNumber:_FillValue = -2147483647 ;
  	string variable_names(nvars) ;
  		string variable_names:_FillValue = "" ;
  data:

   dateTime = -28800, -28800, -28800, -28800, -28800, -28800, -28800, -28800,
      -28800, -28800, -28800, -32400, -32400, -32400, -32400, -32400, -32400,
      -32400, -32400, -32400, -32400, -21600, -21600, -21600, -21600, -21600,
      -21600, -21600, -21600, -21600, -21600, -21600, -21600, -14400, -14400,
      -14400, -14400, -14400, -14400, -14400, -14400, -14400, -14400, 7200,
      7200, 7200, 7200, 7200, 7200, 7200, 7200, 7200, 7200, 7200, 14400,
      14400, 14400, 14400, 14400, 14400, 14400, 14400, 14400, 10800, 10800,
      10800, 10800, 10800, 10800, 10800, 10800, 10800, 3600, 3600, 3600,
      3600, 3600, 3600, 3600, 3600, 3600, 3600, 3600, 3600, 18000, 18000,
      18000, 18000, 18000, 18000, 18000, 18000, 18000, 18000, 18000, 18000,
      18000, 18000, 18000, 18000, 18000, 18000, 18000, 18000, 18000, 3600,
      3600, 3600, 3600, 3600, 3600, 3600, 3600, 3600, 3600, 7200, 7200, 7200,
      7200, 7200, 7200, 7200, 7200, 7200, 7200, 7200, 7200, 7200, 28800,
      28800, 28800, 28800, 28800, 28800, 28800, 28800, 28800, 28800, 28800,
      28800, 28800, 28800, 28800, 28800, 28800, 28800, 28800, 28800, 25200,
      25200, 25200, 25200, 25200, 25200, 25200, 25200, 25200, 25200, 32400,
      32400, 32400, 32400, 32400, 32400, 32400, 32400, 32400, 32400, 32400,
      39600, 39600, 39600, 39600, 39600, 39600, 39600, 39600, 39600, 39600,
      39600, 39600, 39600, 39600, 39600, 39600, 39600, 39600, 39600, 39600,
      39600, 39600, 39600, 36000, 36000, 36000, 36000, 36000, 36000, 36000,
      36000, 36000, 36000, 36000, 36000, 36000, 36000, 36000, 36000, 36000,
      36000, 36000, 36000, 36000, 36000, 36000, 36000, 36000, 36000 ;

   depth = 60, 500, 40, 100, 180, 80, 1, 140, 120, 300, 20, 125, 250, 25,
      150, 200, 1, 300, 50, 500, 75, 10, 300, 140, 120, 500, 100, 80, 180,
      60, 40, 20, 1, 100, 120, 140, 180, 20, 500, 40, 60, 300, 80, 40, 500,
      60, 180, 20, 120, 140, 1, 80, 300, 100, 25, 100, 50, 1, 300, 250, 500,
      125, 200, 75, 25, 500, 250, 150, 300, 50, 200, 100, 100, 180, 300, 40,
      60, 10, 20, 1, 120, 140, 500, 80, 500, 150, 300, 250, 125, 75, 100, 50,
      200, 25, 100, 50, 125, 75, 300, 250, 500, 25, 200, 150, 1, 100, 200,
      50, 1.5, 125, 75, 300, 25, 150, 250, 140, 80, 500, 300, 1, 100, 40, 60,
      10, 20, 180, 5, 120, 300, 140, 1, 120, 100, 80, 500, 40, 180, 60, 80,
      100, 300, 120, 500, 140, 20, 1, 180, 40, 100, 50, 200, 1.5, 125, 75,
      150, 300, 25, 250, 500, 40, 100, 80, 140, 120, 1, 20, 300, 180, 60,
      100, 80, 1, 140, 300, 120, 20, 500, 60, 180, 300, 100, 120, 500, 25,
      140, 20, 5, 40, 180, 60, 45, 80, 60, 300, 80, 4, 1, 120, 5, 140, 100,
      10, 20, 180, 40, 500, 60, 300, 80, 100, 1, 120, 140, 180, 500, 10, 20, 40 ;

   latitude = 8.1, 8.1, 8.1, 8.1, 8.1, 8.1, 8.1, 8.1, 8.1, 8.1, 8.1, -8, -8,
      -8, -8, -8, -8, -8, -8, -8, -8, -4.03686, -4.03686, -4.03686, -4.03686,
      -4.03686, -4.03686, -4.03686, -4.03686, -4.03686, -4.03686, -4.03686,
      -4.03686, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, -5, -5, -5, -5, -5, -5, -5, -5,
      -5, -5, -5, 2, 2, 2, 2, 2, 2, 2, 2, 2, -5, -5, -5, -5, -5, -5, -5, -5,
      -5, -8.01557, -8.01557, -8.01557, -8.01557, -8.01557, -8.01557,
      -8.01557, -8.01557, -8.01557, -8.01557, -8.01557, -8.01557, -2, -2, -2,
      -2, -2, -2, -2, -2, -2, -2, -2.2, -2.2, -2.2, -2.2, -2.2, -2.2, -2.2,
      -2.2, -2.2, -2.2, -2.2, -0.0141, -0.0141, -0.0141, -0.0141, -0.0141,
      -0.0141, -0.0141, -0.0141, -0.0141, -0.0141, 0.00453, 0.00453, 0.00453,
      0.00453, 0.00453, 0.00453, 0.00453, 0.00453, 0.00453, 0.00453, 0.00453,
      0.00453, 0.00453, 2, 2, 2, 2, 2, 2, 2, 2, 2, -8, -8, -8, -8, -8, -8,
      -8, -8, -8, -8, -8, -0.01599, -0.01599, -0.01599, -0.01599, -0.01599,
      -0.01599, -0.01599, -0.01599, -0.01599, -0.01599, 2, 2, 2, 2, 2, 2, 2,
      2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
      0, 0, 0, -6.0014, -6.0014, -6.0014, -6.0014, -6.0014, -6.0014, -6.0014,
      -6.0014, -6.0014, -6.0014, -6.0014, -6.0014, -6.0014, -6.0014,
      -4.03584, -4.03584, -4.03584, -4.03584, -4.03584, -4.03584, -4.03584,
      -4.03584, -4.03584, -4.03584, -4.03584, -4.03584 ;

   longitude = -125, -125, -125, -125, -125, -125, -125, -125, -125, -125,
      -125, 164.8, 164.8, 164.8, 164.8, 164.8, 164.8, 164.8, 164.8, 164.8,
      164.8, 67.24096, 67.24096, 67.24096, 67.24096, 67.24096, 67.24096,
      67.24096, 67.24096, 67.24096, 67.24096, 67.24096, 67.24096, -140, -140,
      -140, -140, -140, -140, -140, -140, -140, -140, -139.9, -139.9, -139.9,
      -139.9, -139.9, -139.9, -139.9, -139.9, -139.9, -139.9, -139.9, 165.2,
      165.2, 165.2, 165.2, 165.2, 165.2, 165.2, 165.2, 165.2, 165.2, 165.2,
      165.2, 165.2, 165.2, 165.2, 165.2, 165.2, 165.2, 80.45833, 80.45833,
      80.45833, 80.45833, 80.45833, 80.45833, 80.45833, 80.45833, 80.45833,
      80.45833, 80.45833, 80.45833, -155, -155, -155, -155, -155, -155, -155,
      -155, -155, -155, -170, -170, -170, -170, -170, -170, -170, -170, -170,
      -170, -170, 155.9603, 155.9603, 155.9603, 155.9603, 155.9603, 155.9603,
      155.9603, 155.9603, 155.9603, 155.9603, -22.98389, -22.98389,
      -22.98389, -22.98389, -22.98389, -22.98389, -22.98389, -22.98389,
      -22.98389, -22.98389, -22.98389, -22.98389, -22.98389, -110, -110,
      -110, -110, -110, -110, -110, -110, -110, -110.1, -110.1, -110.1,
      -110.1, -110.1, -110.1, -110.1, -110.1, -110.1, -110.1, -110.1,
      155.957, 155.957, 155.957, 155.957, 155.957, 155.957, 155.957, 155.957,
      155.957, 155.957, -140, -140, -140, -140, -140, -140, -140, -140, -140,
      -140, -140, -125.1, -125.1, -125.1, -125.1, -125.1, -125.1, -125.1,
      -125.1, -125.1, -125.1, -139.9, -139.9, -139.9, -139.9, -139.9, -139.9,
      -139.9, -139.9, -139.9, -139.9, -139.9, -139.9, -139.9, 8.00453,
      8.00453, 8.00453, 8.00453, 8.00453, 8.00453, 8.00453, 8.00453, 8.00453,
      8.00453, 8.00453, 8.00453, 8.00453, 8.00453, 67.242, 67.242, 67.242,
      67.242, 67.242, 67.242, 67.242, 67.242, 67.242, 67.242, 67.242, 67.242 ;

   sequenceNumber = 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 2, 2, 2, 2, 2, 2, 2, 2,
      2, 2, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4,
      5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 6, 6, 6, 6, 6, 6, 6, 6, 6, 7, 7, 7, 7,
      7, 7, 7, 7, 7, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9,
      9, 9, 9, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 11, 11, 11, 11,
      11, 11, 11, 11, 11, 11, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12,
      12, 13, 13, 13, 13, 13, 13, 13, 13, 13, 14, 14, 14, 14, 14, 14, 14, 14,
      14, 14, 14, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 16, 16, 16, 16, 16,
      16, 16, 16, 16, 16, 16, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 18, 18,
      18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 19, 19, 19, 19, 19, 19, 19,
      19, 19, 19, 19, 19, 19, 19, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20 ;

   variable_names = "sea_water_salinity", "sea_water_temperature" ;
  } // group MetaData

group: ObsError {
  variables:
  	float salinity(Location) ;
  		salinity:_FillValue = 9.96921e+36f ;
  	float waterTemperature(Location) ;
  		waterTemperature:_FillValue = 9.96921e+36f ;
  data:

   salinity = 0.2522745, 0.1063194, 0.2849693, 0.166195, 0.09365788,
      0.200834, 0.2371611, 0.08366414, 0.1299536, 0.1010965, 0.1687779,
      0.7850429, 0.4356464, 1.591666, 0.8089812, 0.6832849, 1.697105,
      0.3133486, 1.511612, 0.2497392, 1.203681, 0.2197831, 0.1222905,
      0.08824342, 0.1645312, 0.1172962, 0.1364866, 0.1435371, 0.1202509,
      0.2682254, 0.1998587, 0.1259456, 0.6451571, 1.210507, 1.097976,
      0.8719119, 0.4586407, 1.158771, 0.1140179, 1.141717, 1.164443,
      0.1429435, 1.197306, 0.2177143, 0.1228545, 0.2259728, 0.1939958,
      0.2478939, 0.2443465, 0.2529505, 0.3637651, 0.2088105, 0.1383288,
      0.1579156, 0.1400251, 0.27416, 0.2761041, 0.2834496, 0.1044707,
      0.1786518, 0.117582, 0.1529245, 0.224429, 1.179957, 1.548487,
      0.2490613, 0.510761, 0.9821573, 0.3357151, 1.441269, 0.880218, 0.92051,
      0.1224098, 0.0733786, 0.09151919, 0.3130135, 0.3720615, 0.1560941,
      0.1031811, 0.2011424, 0.2196218, 0.06576524, 0.09795111, 0.1263566,
      0.1404088, 1.438963, 0.1937371, 0.2689984, 1.490757, 1.047074,
      1.288639, 1.00524, 0.6400538, 1.021853, 0.1832772, 0.181006, 0.1896285,
      0.2019524, 0.1270845, 0.2043958, 0.1171445, 0.2605884, 0.2675938,
      0.2263254, 0.3653024, 0.2850498, 0.2288099, 0.09864562, 0.1805917,
      0.3270485, 0.1413604, 0.1385984, 0.215419, 0.1264153, 0.1776507,
      0.2440303, 0.391326, 0.174588, 0.1708031, 0.05932364, 0.3705409,
      0.2244651, 0.1368625, 0.1493623, 0.05727173, 0.166375, 0.05866817,
      0.2646765, 0.1636383, 0.6282568, 1.789018, 0.735101, 0.8842987,
      1.167529, 0.1027457, 1.507743, 0.4915881, 1.568499, 1.363651, 1.080779,
      0.1952056, 0.9173244, 0.06207152, 0.757747, 1.901986, 1.914773,
      0.5039916, 1.71778, 0.2737243, 0.09864481, 0.2359564, 0.3332464,
      0.3405225, 0.1123013, 0.1469922, 0.0873469, 0.2929741, 0.1750725,
      0.1346339, 0.138216, 0.2096565, 0.1308088, 0.1126329, 0.2334442,
      0.2602245, 0.1921947, 0.1253058, 0.09266749, 0.155894, 0.1143336,
      0.1697396, 0.2593261, 0.1232226, 0.1157582, 0.1466153, 0.1364038,
      0.1281689, 0.2194774, 0.09342678, 0.1313902, 0.05775158, 0.09673796,
      0.1344558, 0.3084517, 0.2484634, 0.3372627, 0.3816409, 0.1399285,
      0.1459216, 0.2595628, 0.151517, 0.2104556, 0.1805469, 0.1823283,
      0.2343753, 1.871043, 1.056106, 0.1652864, 1.759668, 0.2059344,
      0.1846005, 0.8090061, 0.5420793, 0.1961852, 0.1148487, 0.1676946,
      0.1995637, 0.1171088, 0.2132636, 0.1414041, 0.6741951, 0.2209578,
      0.06775443, 0.1180433, 0.1100427, 0.2316091, 0.2603508, 0.1870268 ;

   waterTemperature = 1.743426, 0.5193261, 1.494207, 0.8796794, 0.5286709,
      1.343593, 0.5824349, 0.61001, 0.667032, 0.5093725, 0.8844231,
      0.9340492, 1.007331, 0.468168, 0.9813886, 1.036275, 0.5447601,
      0.770175, 0.3583136, 0.6713341, 0.8158218, 0.7916454, 0.6055509,
      0.7106637, 0.7956954, 0.5452055, 1.114186, 1.488101, 0.6829131,
      1.468622, 1.12228, 0.7781153, 0.9701674, 1.599963, 1.476451, 0.7450125,
      0.5824413, 0.644627, 0.6039046, 0.8115129, 0.903461, 0.5930381,
      1.065919, 0.2801136, 0.5537068, 0.737125, 0.8197537, 0.3324322,
      1.362025, 1.135762, 0.3594703, 1.020024, 0.6098969, 1.323719,
      0.4565539, 0.5973899, 0.5753483, 0.272785, 0.5647165, 0.9110706,
      0.5528083, 1.167597, 1.235241, 0.5491017, 0.4130876, 0.589695,
      1.195557, 0.9150438, 0.7125937, 0.4867784, 1.229869, 0.6954335,
      0.9935142, 0.6311837, 0.5309837, 1.439539, 1.658565, 0.6073291,
      0.5337266, 0.7063531, 0.8778601, 0.7684838, 0.4986047, 1.235635,
      0.5999914, 1.308395, 0.5793702, 0.7610333, 0.9590447, 0.6941347,
      0.7923799, 0.4928668, 1.169785, 0.2800499, 0.7219963, 0.3700807,
      0.8848718, 0.4830801, 0.5760365, 0.8778846, 0.5401599, 0.3846734,
      1.235485, 1.295008, 0.3513189, 0.466359, 1.139407, 0.4031729,
      0.5074973, 1.204991, 0.4061031, 0.6839842, 0.4782485, 1.380711,
      0.8387715, 0.7210994, 1.324711, 0.6442875, 0.6358635, 1.226067,
      1.129524, 1.05598, 1.353591, 0.5635409, 0.6810182, 0.6161842,
      0.9409899, 0.9163142, 0.5753275, 0.5561668, 1.119911, 0.5457644,
      0.6782846, 1.336049, 0.5781834, 1.43989, 0.5525411, 1.019478, 1.248575,
      1.2796, 0.5426413, 1.302236, 0.5345117, 1.036997, 0.6088989, 0.4321637,
      0.6309587, 0.7555988, 0.4618859, 0.403173, 1.153354, 0.3227628,
      1.173669, 0.4006487, 1.37786, 0.6794108, 0.3855352, 0.8370423,
      0.6134599, 0.7724864, 1.520247, 1.046432, 0.8824214, 1.474335,
      0.5206715, 0.4941791, 0.5990528, 0.5935799, 0.8832166, 1.424629,
      1.542141, 0.8646343, 0.6747602, 0.5828347, 0.8573534, 0.8243105,
      0.5863172, 1.030508, 0.5895203, 0.6056085, 1.342003, 1.028111,
      0.6016723, 0.527028, 1.005599, 0.5325223, 0.5584281, 0.5712408,
      0.7219398, 0.8380678, 0.6462824, 1.317487, 0.8282857, 0.6612134,
      0.7838165, 1.337059, 1.043711, 0.6533467, 1.208123, 0.638188,
      0.6995534, 1.724898, 1.705356, 0.6825911, 1.242171, 0.6282559, 1.50075,
      0.5917126, 1.514512, 1.116175, 0.5734112, 0.8052191, 0.656361,
      0.668393, 0.5316752, 0.5864132, 0.8440492, 1.121295 ;
  } // group ObsError

group: ObsValue {
  variables:
  	float salinity(Location) ;
  		salinity:_FillValue = 9.96921e+36f ;
  	float waterTemperature(Location) ;
  		waterTemperature:_FillValue = 9.96921e+36f ;
  data:

   salinity = 34.57398, 34.60444, 34.41549, 34.71024, 34.73309, 34.662,
      34.34, 34.74724, 34.74189, 34.7036, 34.24408, 35.5955, 35.39627,
      34.81105, 35.6922, 35.70549, 34.74729, 35.04684, 34.93018, 34.64479,
      35.09085, 35.47, 35.0326, 35.15076, 35.16211, 34.8932, 35.23, 35.20581,
      35.15009, 35.18, 35.49, 35.05608, 34.98, 35.07314, 34.85984, 34.85921,
      34.88235, 34.99768, 34.61454, 35.01868, 35.04686, 34.82505, 35.07153,
      35.2707, 34.63697, 35.37906, 35.02031, 35.21252, 35.3908, 35.29946,
      35.5, 35.45095, 34.8038, 35.52097, 34.64267, 35.20449, 34.78244, 34.83,
      34.80511, 34.77232, 34.66197, 35.34407, 35.05775, 35.1338, 34.75198,
      34.61681, 35.2095, 35.6226, 34.84489, 34.90092, 35.87683, 35.35735,
      34.69, 34.86082, 34.85189, 34.26, 34.66, 34.25, 34.25, 34.22, 34.85972,
      34.86072, 34.7815, 34.88726, 34.59576, 35.50129, 34.79575, 34.79715,
      35.4471, 35.26348, 35.33844, 35.21389, 35.02264, 35.18464, 35.43448,
      35.26216, 35.48049, 35.34953, 34.76404, 34.85212, 34.62323, 35.22366,
      35.13306, 35.57404, 35.59, 34.81, 35.11, 34.76, 34.58, 35.05, 34.64,
      34.87, 34.63, 35.4, 34.93, 35.50653, 36.38, 34.69085, 35.17369, 36.34,
      35.78912, 36.34, 36.5, 36.34, 36.32, 35.40076, 36.34, 35.75, 34.83435,
      34.89127, 33.98383, 34.91024, 34.93637, 34.95012, 34.65226, 34.64199,
      34.87164, 35.51104, 35.61652, 35.54525, 34.79385, 35.31134, 34.66566,
      34.98342, 35.08948, 34.9439, 34.86064, 35.28613, 34.75, 34.77, 35.11,
      34.36, 35.01, 34.64, 35.4, 34.88, 34.63, 34.89, 34.61314, 35.01323,
      35.08269, 35.07761, 34.87947, 34.9267, 35.13, 35.0029, 34.83858,
      34.89431, 35.04663, 34.93151, 34.92387, 34.79, 34.87672, 34.83274,
      34.90145, 34.66761, 34.63993, 34.84803, 34.85432, 34.86982, 35.09964,
      35.33, 34.64524, 35.07434, 35.08952, 35.07367, 35.33, 35.28, 34.97347,
      35.25, 35.0976, 35.33, 35.93, 35.11495, 35.88, 32.29442, 32.71, 35.77,
      34.71, 35.64164, 35.72212, 34.94, 35.95, 35.54502, 35.98, 34.68404,
      35.16, 35.02942, 35.19083, 35.32, 34.97, 35.14178, 35.14002, 35.13965,
      34.91897, 35.51, 35.05788, 35.32 ;

   waterTemperature = 18.94, 8.149994, 25.89001, 12.94, 11.30002, 14.42001,
      28.22, 12.01001, 12.39001, 10.25, 27.92999, 26.25, 17.27002, 29.42001,
      25.02002, 21.20999, 29.70999, 13.76001, 29.39999, 8.540009, 29.45999,
      29.97, 11.80002, 15.84, 16.70999, 9.220001, 17.36002, 20.63, 15.09,
      25.67999, 28.75, 29.85001, 30.67001, 21.70999, 14.85001, 13.86002,
      13.03, 26.5, 7.730011, 26.08002, 24.77002, 11.39999, 23.86002,
      27.74002, 8.110016, 27.74002, 14.10001, 27.74002, 20.34, 17.99002,
      27.72, 26.47, 10.87, 24.57001, 29.87, 28.78, 29.60001, 29.87, 11.45999,
      12.24002, 8.779999, 28.67001, 17.91, 29.57001, 29.92001, 8.070007,
      15.52002, 27.69, 11.47, 29.84, 24.01001, 29.29001, 15.58002, 12.26001,
      10.45001, 28.35001, 20.79001, 28.64999, 28.58002, 28.92001, 14.34,
      13.54001, 8.660004, 17.22, 7.52002, 23.42999, 11.08002, 11.32001,
      25.39001, 27.10001, 26.20001, 27.45001, 14.85001, 27.45001, 28.13,
      28.47, 26.83002, 28.33002, 10.67999, 12.14001, 8.300018, 28.39999,
      16.5, 25.70999, 28.38, 29.67999, 16.94, 29.79001, 30.12, 29.62, 29.78,
      12.27002, 29.91, 23.85001, 13.63, 15.27002, 20.57001, 7.630005,
      12.20001, 28.36002, 17.80002, 26.94, 24.04001, 27.72, 27.58002, 14.34,
      27.78, 16.24002, 11.86002, 13.97, 28.62, 14.23001, 14.45001, 15.23001,
      8.670013, 24.42999, 13.44, 25.57001, 23.22, 20.17001, 10.92001, 17.47,
      8.589996, 14.11002, 26.91, 26.99002, 12.51001, 26.29001, 29.70001,
      29.80002, 17.02002, 29.89999, 29.63, 29.78, 24.29001, 12.38, 29.91,
      13.70999, 7.700012, 26.26001, 22.04001, 24.19, 14.22, 16.35001,
      26.54001, 26.41, 11.58002, 13.20001, 24.92999, 16.39999, 22.87,
      27.77002, 14.32001, 11.64999, 15, 26.77002, 8.360016, 25.16, 13.47,
      11.99002, 19.89999, 18.64001, 8.330017, 26.28, 16.95999, 26.29001,
      26.45999, 26.12, 14.08002, 25.75, 26.05002, 24.57001, 18.53, 11.66,
      17.61002, 29.07001, 29.34, 16.47, 28.64999, 16.02002, 16.95001, 28.28,
      23.87, 15.17001, 19.38, 7.420013, 25.79001, 11.75, 19.97, 17.08002,
      30.25, 16.03, 15.5, 14.81, 9.410004, 30.12, 29.95001, 28.56 ;
  } // group ObsValue

group: PreQC {
  variables:
  	float salinity(Location) ;
  		salinity:_FillValue = 9.96921e+36f ;
  	float waterTemperature(Location) ;
  		waterTemperature:_FillValue = 9.96921e+36f ;
  data:

   salinity = 0.08789432, 0.08789432, 0.08789432, 0.08789432, 0.08789432,
      0.08789432, 0.08789432, 0.08789432, 0.08789432, 0.08789432, 0.08789432,
      0.2789434, 0.2789434, 0.2789434, 0.2789434, 0.2789434, 0.2789434,
      0.2789434, 0.2789434, 0.2789434, 0.2789434, 0.4881761, 0.4881761,
      0.4881761, 0.4881761, 0.4881761, 0.4881761, 0.4881761, 0.4881761,
      0.4881761, 0.4881761, 0.4881761, 0.4881761, 0.09344757, 0.09344757,
      0.09344757, 0.09344757, 0.09344757, 0.09344757, 0.09344757, 0.09344757,
      0.09344757, 0.09344757, 0.3562652, 0.3562652, 0.3562652, 0.3562652,
      0.3562652, 0.3562652, 0.3562652, 0.3562652, 0.3562652, 0.3562652,
      0.3562652, 0.6465657, 0.6465657, 0.6465657, 0.6465657, 0.6465657,
      0.6465657, 0.6465657, 0.6465657, 0.6465657, 0.245206, 0.245206,
      0.245206, 0.245206, 0.245206, 0.245206, 0.245206, 0.245206, 0.245206,
      0.344362, 0.344362, 0.344362, 0.344362, 0.344362, 0.344362, 0.344362,
      0.344362, 0.344362, 0.344362, 0.344362, 0.344362, 0.2459739, 0.2459739,
      0.2459739, 0.2459739, 0.2459739, 0.2459739, 0.2459739, 0.2459739,
      0.2459739, 0.2459739, 0.2994778, 0.2994778, 0.2994778, 0.2994778,
      0.2994778, 0.2994778, 0.2994778, 0.2994778, 0.2994778, 0.2994778,
      0.2994778, 0.3914765, 0.3914765, 0.3914765, 0.3914765, 0.3914765,
      0.3914765, 0.3914765, 0.3914765, 0.3914765, 0.3914765, 0.6239262,
      0.6239262, 0.6239262, 0.6239262, 0.6239262, 0.6239262, 0.6239262,
      0.6239262, 0.6239262, 0.6239262, 0.6239262, 0.6239262, 0.6239262,
      0.1783193, 0.1783193, 0.1783193, 0.1783193, 0.1783193, 0.1783193,
      0.1783193, 0.1783193, 0.1783193, 0.1653826, 0.1653826, 0.1653826,
      0.1653826, 0.1653826, 0.1653826, 0.1653826, 0.1653826, 0.1653826,
      0.1653826, 0.1653826, 0.5274251, 0.5274251, 0.5274251, 0.5274251,
      0.5274251, 0.5274251, 0.5274251, 0.5274251, 0.5274251, 0.5274251,
      0.3551692, 0.3551692, 0.3551692, 0.3551692, 0.3551692, 0.3551692,
      0.3551692, 0.3551692, 0.3551692, 0.3551692, 0.3551692, 0.2711022,
      0.2711022, 0.2711022, 0.2711022, 0.2711022, 0.2711022, 0.2711022,
      0.2711022, 0.2711022, 0.2711022, 0.4063673, 0.4063673, 0.4063673,
      0.4063673, 0.4063673, 0.4063673, 0.4063673, 0.4063673, 0.4063673,
      0.4063673, 0.4063673, 0.4063673, 0.4063673, 0.3125914, 0.3125914,
      0.3125914, 0.3125914, 0.3125914, 0.3125914, 0.3125914, 0.3125914,
      0.3125914, 0.3125914, 0.3125914, 0.3125914, 0.3125914, 0.3125914,
      0.4828305, 0.4828305, 0.4828305, 0.4828305, 0.4828305, 0.4828305,
      0.4828305, 0.4828305, 0.4828305, 0.4828305, 0.4828305, 0.4828305 ;

   waterTemperature = 0.3304284, 0.3304284, 0.3304284, 0.3304284, 0.3304284,
      0.3304284, 0.3304284, 0.3304284, 0.3304284, 0.3304284, 0.3304284,
      0.4522219, 0.4522219, 0.4522219, 0.4522219, 0.4522219, 0.4522219,
      0.4522219, 0.4522219, 0.4522219, 0.4522219, 0.5740165, 0.5740165,
      0.5740165, 0.5740165, 0.5740165, 0.5740165, 0.5740165, 0.5740165,
      0.5740165, 0.5740165, 0.5740165, 0.5740165, 0.3443506, 0.3443506,
      0.3443506, 0.3443506, 0.3443506, 0.3443506, 0.3443506, 0.3443506,
      0.3443506, 0.3443506, 0.2669469, 0.2669469, 0.2669469, 0.2669469,
      0.2669469, 0.2669469, 0.2669469, 0.2669469, 0.2669469, 0.2669469,
      0.2669469, 0.5118217, 0.5118217, 0.5118217, 0.5118217, 0.5118217,
      0.5118217, 0.5118217, 0.5118217, 0.5118217, 0.4708711, 0.4708711,
      0.4708711, 0.4708711, 0.4708711, 0.4708711, 0.4708711, 0.4708711,
      0.4708711, 0.3297694, 0.3297694, 0.3297694, 0.3297694, 0.3297694,
      0.3297694, 0.3297694, 0.3297694, 0.3297694, 0.3297694, 0.3297694,
      0.3297694, 0.7652588, 0.7652588, 0.7652588, 0.7652588, 0.7652588,
      0.7652588, 0.7652588, 0.7652588, 0.7652588, 0.7652588, 0.399832,
      0.399832, 0.399832, 0.399832, 0.399832, 0.399832, 0.399832, 0.399832,
      0.399832, 0.399832, 0.399832, 0.4094992, 0.4094992, 0.4094992,
      0.4094992, 0.4094992, 0.4094992, 0.4094992, 0.4094992, 0.4094992,
      0.4094992, 0.7739636, 0.7739636, 0.7739636, 0.7739636, 0.7739636,
      0.7739636, 0.7739636, 0.7739636, 0.7739636, 0.7739636, 0.7739636,
      0.7739636, 0.7739636, 0.5043824, 0.5043824, 0.5043824, 0.5043824,
      0.5043824, 0.5043824, 0.5043824, 0.5043824, 0.5043824, 0.4389331,
      0.4389331, 0.4389331, 0.4389331, 0.4389331, 0.4389331, 0.4389331,
      0.4389331, 0.4389331, 0.4389331, 0.4389331, 0.3698398, 0.3698398,
      0.3698398, 0.3698398, 0.3698398, 0.3698398, 0.3698398, 0.3698398,
      0.3698398, 0.3698398, 0.2308534, 0.2308534, 0.2308534, 0.2308534,
      0.2308534, 0.2308534, 0.2308534, 0.2308534, 0.2308534, 0.2308534,
      0.2308534, 0.5125766, 0.5125766, 0.5125766, 0.5125766, 0.5125766,
      0.5125766, 0.5125766, 0.5125766, 0.5125766, 0.5125766, 0.3485442,
      0.3485442, 0.3485442, 0.3485442, 0.3485442, 0.3485442, 0.3485442,
      0.3485442, 0.3485442, 0.3485442, 0.3485442, 0.3485442, 0.3485442,
      0.3094093, 0.3094093, 0.3094093, 0.3094093, 0.3094093, 0.3094093,
      0.3094093, 0.3094093, 0.3094093, 0.3094093, 0.3094093, 0.3094093,
      0.3094093, 0.3094093, 0.5460482, 0.5460482, 0.5460482, 0.5460482,
      0.5460482, 0.5460482, 0.5460482, 0.5460482, 0.5460482, 0.5460482,
      0.5460482, 0.5460482 ;
  } // group PreQC
}
