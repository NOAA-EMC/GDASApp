netcdf rads_adt_c2_2018104.tmp {
dimensions:
	time = UNLIMITED ; // (11 currently)
variables:
	int adt_egm2008(time) ;
		adt_egm2008:_FillValue = 2147483647 ;
		adt_egm2008:long_name = "absolute dynamic topography (EGM2008)" ;
		adt_egm2008:standard_name = "absolute_dynamic_topography_egm2008" ;
		adt_egm2008:units = "m" ;
		adt_egm2008:scale_factor = 0.0001 ;
		adt_egm2008:coordinates = "lon lat" ;
	int adt_xgm2016(time) ;
		adt_xgm2016:_FillValue = 2147483647 ;
		adt_xgm2016:long_name = "absolute dynamic topography (XGM2016)" ;
		adt_xgm2016:standard_name = "absolute_dynamic_topography_xgm2016" ;
		adt_xgm2016:units = "m" ;
		adt_xgm2016:scale_factor = 0.0001 ;
		adt_xgm2016:coordinates = "lon lat" ;
	int cycle(time) ;
		cycle:_FillValue = 2147483647 ;
		cycle:long_name = "cycle number" ;
		cycle:field = 9905s ;
	int lat(time) ;
		lat:_FillValue = 2147483647 ;
		lat:long_name = "latitude" ;
		lat:standard_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:scale_factor = 1.e-07 ;
		lat:field = 201s ;
		lat:comment = "Positive latitude is North latitude, negative latitude is South latitude" ;
	int lon(time) ;
		lon:_FillValue = 2147483647 ;
		lon:long_name = "longitude" ;
		lon:standard_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:scale_factor = 1.e-07 ;
		lon:field = 301s ;
		lon:comment = "East longitude relative to Greenwich meridian" ;
	int pass(time) ;
		pass:_FillValue = 2147483647 ;
		pass:long_name = "pass number" ;
		pass:field = 9906s ;
	short sla(time) ;
		sla:_FillValue = 32767s ;
		sla:long_name = "sea level anomaly" ;
		sla:standard_name = "sea_surface_height_above_sea_level" ;
		sla:units = "m" ;
		sla:quality_flag = "swh sig0 range_rms range_numval flags peakiness" ;
		sla:scale_factor = 0.0001 ;
		sla:coordinates = "lon lat" ;
		sla:field = 0s ;
		sla:comment = "Sea level determined from satellite altitude - range - all altimetric corrections" ;
	double time_mjd(time) ;
		time_mjd:long_name = "Modified Julian Days" ;
		time_mjd:standard_name = "time" ;
		time_mjd:units = "days since 1858-11-17 00:00:00 UTC" ;
		time_mjd:field = 105s ;
		time_mjd:comment = "UTC time of measurement expressed in Modified Julian Days" ;

// global attributes:
		:Conventions = "CF-1.7" ;
		:title = "RADS 4 pass file" ;
		:institution = "EUMETSAT / NOAA / TU Delft" ;
		:source = "radar altimeter" ;
		:references = "RADS Data Manual, Version 4.2 or later" ;
		:featureType = "trajectory" ;
		:ellipsoid = "TOPEX" ;
		:ellipsoid_axis = 6378136.3 ;
		:ellipsoid_flattening = 0.00335281317789691 ;
		:filename = "rads_adt_c2_2018104.nc" ;
		:mission_name = "CRYOSAT2" ;
		:mission_phase = "a" ;
		:log01 = "2019-01-11 | rads2nc --ymd=180414000000,180415000000 -C1,1000 -Sc2 -Vadt_egm2008,adt_xgm2016,sla,time_mjd,lon,lat,cycle,pass -Xxgm2016 -Xadt.xml -o/ftp/rads/adt//2018/rads_adt_c2_2018104.nc: RAW data from" ;
		:history = "Fri Jan 26 15:44:21 2024: ncks -d time,0,10 /scratch1/NCEPDEV/stmp4/Shastri.Paturi/forAndrew/gdas.20180414/00/adt/rads_adt_c2_2018104.nc rads_adt_c2_2018104.tmp.nc\n",
			"2019-01-11 12:29:35 : rads2nc --ymd=180414000000,180415000000 -C1,1000 -Sc2 -Vadt_egm2008,adt_xgm2016,sla,time_mjd,lon,lat,cycle,pass -Xxgm2016 -Xadt.xml -o/ftp/rads/adt//2018/rads_adt_c2_2018104.nc" ;
		:NCO = "netCDF Operators version 5.0.6 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco)" ;
data:

 adt_egm2008 = 11661, 11735, 12134, 11616, 12174, 11993, 12093, 11915, 11687, 
    10992, 11465 ;

 adt_xgm2016 = 11996, 12167, 12391, 11456, 11614, 11219, 11324, 11333, 11465, 
    11170, 11951 ;

 cycle = 104, 104, 104, 104, 104, 104, 104, 104, 104, 104, 104 ;

 lat = -251089129, -250517057, -249944976, -249372888, -248800790, 
    -248228689, -247656580, -247084459, -246512330, -245940194, -245368050 ;

 lon = 738495892, 738432015, 738368162, 738304331, 738240522, 738176735, 
    738112971, 738049229, 737985509, 737921811, 737858134 ;

 pass = 285, 285, 285, 285, 285, 285, 285, 285, 285, 285, 285 ;

 sla = 2359, 2193, 2585, 2183, 2651, 2317, 2454, 2384, 2214, 1494, 1956 ;

 time_mjd = 58222.0000010569, 58222.0000119763, 58222.0000228957, 
    58222.0000338151, 58222.0000447346, 58222.0000556539, 58222.0000665733, 
    58222.0000774927, 58222.0000884121, 58222.0000993315, 58222.0001102509 ;
}
