netcdf output_2 {
dimensions:
	Scanline = 6 ;
	Field_of_view = 5 ;
	Channel = 22 ;
	Qc_dim = 4 ;
variables:
	short Atm_type(Scanline, Field_of_view) ;
		Atm_type:description = "type of atmosphere:currently missing" ;
		Atm_type:coordinates = "Longitude Latitude" ;
	short BT(Scanline, Field_of_view, Channel) ;
		BT:long_name = "Channel Temperature (K)" ;
		BT:units = "Kelvin" ;
		BT:coordinates = "Longitude Latitude Freq" ;
		BT:scale_factor = 0.01 ;
		BT:_FillValue = -999s ;
		BT:valid_range = 0, 50000 ;
	short CLW(Scanline, Field_of_view) ;
		CLW:long_name = "Cloud liquid Water (mm)" ;
		CLW:units = "mm" ;
		CLW:coordinates = "Longitude Latitude" ;
		CLW:scale_factor = 0.01 ;
		CLW:_FillValue = -999s ;
		CLW:valid_range = 0, 10000 ;
	short ChanSel(Scanline, Field_of_view, Channel) ;
		ChanSel:long_name = "Channels Selection Used in Retrieval" ;
		ChanSel:units = "1" ;
		ChanSel:coordinates = "Longitude Latitude Freq" ;
		ChanSel:_FillValue = -999s ;
		ChanSel:valid_range = 0, 1 ;
	float ChiSqr(Scanline, Field_of_view) ;
		ChiSqr:description = "Convergence rate: <3-good,>10-bad" ;
		ChiSqr:units = "1" ;
		ChiSqr:coordinates = "Longitude Latitude" ;
		ChiSqr:_FillValue = -999.f ;
		ChiSqr:valid_range = 0.f, 1000.f ;
	short CldBase(Scanline, Field_of_view) ;
		CldBase:long_name = "Cloud Base Pressure" ;
		CldBase:scale_factor = 0.1 ;
		CldBase:coordinates = "Longitude Latitude" ;
	short CldThick(Scanline, Field_of_view) ;
		CldThick:long_name = "Cloud Thickness" ;
		CldThick:scale_factor = 0.1 ;
		CldThick:coordinates = "Longitude Latitude" ;
	short CldTop(Scanline, Field_of_view) ;
		CldTop:long_name = "Cloud Top Pressure" ;
		CldTop:scale_factor = 0.1 ;
		CldTop:coordinates = "Longitude Latitude" ;
	short Emis(Scanline, Field_of_view, Channel) ;
		Emis:long_name = "Channel Emissivity" ;
		Emis:units = "1" ;
		Emis:coordinates = "Longitude Latitude Freq" ;
		Emis:scale_factor = 0.0001 ;
		Emis:_FillValue = -999s ;
		Emis:valid_range = 0, 10000 ;
	float Freq(Channel) ;
		Freq:description = "Central Frequencies (GHz)" ;
	short GWP(Scanline, Field_of_view) ;
		GWP:long_name = "Graupel Water Path (mm)" ;
		GWP:units = "mm" ;
		GWP:coordinates = "Longitude Latitude" ;
		GWP:scale_factor = 0.01 ;
		GWP:_FillValue = -999s ;
		GWP:valid_range = 0, 10000 ;
	short IWP(Scanline, Field_of_view) ;
		IWP:long_name = "Ice Water Path (mm)" ;
		IWP:units = "mm" ;
		IWP:coordinates = "Longitude Latitude" ;
		IWP:scale_factor = 0.01 ;
		IWP:_FillValue = -999s ;
		IWP:valid_range = 0, 10000 ;
	short LWP(Scanline, Field_of_view) ;
		LWP:long_name = "Liquid Water Path (mm)" ;
		LWP:units = "mm" ;
		LWP:coordinates = "Longitude Latitude" ;
		LWP:scale_factor = 0.01 ;
		LWP:_FillValue = -999s ;
		LWP:valid_range = 0, 10000 ;
	float LZ_angle(Scanline, Field_of_view) ;
		LZ_angle:long_name = "Local Zenith Angle degree" ;
		LZ_angle:units = "degrees" ;
		LZ_angle:coordinates = "Longitude Latitude" ;
		LZ_angle:_FillValue = -999.f ;
		LZ_angle:valid_range = -70.f, 70.f ;
	float Latitude(Scanline, Field_of_view) ;
		Latitude:long_name = "Latitude of the view (-90,90)" ;
		Latitude:units = "degrees" ;
		Latitude:_FillValue = -999.f ;
		Latitude:valid_range = -90.f, 90.f ;
	float Longitude(Scanline, Field_of_view) ;
		Longitude:long_name = "Longitude of the view (-180,180)" ;
		Longitude:units = "degrees" ;
		Longitude:_FillValue = -999.f ;
		Longitude:valid_range = -180.f, 180.f ;
	short Orb_mode(Scanline) ;
		Orb_mode:description = "0-ascending,1-descending" ;
		Orb_mode:units = "1" ;
		Orb_mode:_FillValue = -999s ;
		Orb_mode:valid_range = 0, 1 ;
	short Polo(Channel) ;
		Polo:description = "Polarizations" ;
	short PrecipType(Scanline, Field_of_view) ;
		PrecipType:long_name = "Precipitation Type (Frozen/Liquid)" ;
		PrecipType:coordinates = "Longitude Latitude" ;
	short Prob_SF(Scanline, Field_of_view) ;
		Prob_SF:long_name = "Probability of falling snow (%)" ;
		Prob_SF:units = "percent" ;
		Prob_SF:coordinates = "Longitude Latitude" ;
		Prob_SF:_FillValue = -999s ;
		Prob_SF:valid_range = 0, 100 ;
	short Qc(Scanline, Field_of_view, Qc_dim) ;
		Qc:description = "Qc: 0-good, 1-usable with problem, 2-bad" ;
	float RAzi_angle(Scanline, Field_of_view) ;
		RAzi_angle:long_name = "Relative Azimuth Angle 0-360 degree" ;
		RAzi_angle:coordinates = "Longitude Latitude" ;
	short RFlag(Scanline, Field_of_view) ;
		RFlag:long_name = "Rain Flag" ;
		RFlag:coordinates = "Longitude Latitude" ;
	short RR(Scanline, Field_of_view) ;
		RR:long_name = "Rain Rate (mm/hr)" ;
		RR:units = "mm/hr" ;
		RR:coordinates = "Longitude Latitude" ;
		RR:scale_factor = 0.1 ;
		RR:_FillValue = -999s ;
		RR:valid_range = 0, 1000 ;
	short RWP(Scanline, Field_of_view) ;
		RWP:long_name = "Rain Water Path (mm)" ;
		RWP:units = "mm" ;
		RWP:coordinates = "Longitude Latitude" ;
		RWP:scale_factor = 0.01 ;
		RWP:_FillValue = -999s ;
		RWP:valid_range = 0, 10000 ;
	short SFR(Scanline, Field_of_view) ;
		SFR:long_name = "Snow Fall Rate in mm/hr" ;
		SFR:units = "mm/hr" ;
		SFR:coordinates = "Longitude Latitude" ;
		SFR:scale_factor = 0.01 ;
		SFR:_FillValue = -999s ;
		SFR:valid_range = 0, 10000 ;
	short SIce(Scanline, Field_of_view) ;
		SIce:long_name = "Sea Ice Concentration (%)" ;
		SIce:units = "percent" ;
		SIce:coordinates = "Longitude Latitude" ;
		SIce:_FillValue = -999s ;
		SIce:valid_range = 0, 100 ;
	short SIce_FY(Scanline, Field_of_view) ;
		SIce_FY:long_name = "First-Year Sea Ice Concentration (%)" ;
		SIce_FY:units = "percent" ;
		SIce_FY:coordinates = "Longitude Latitude" ;
		SIce_FY:_FillValue = -999s ;
		SIce_FY:valid_range = 0, 100 ;
	short SIce_MY(Scanline, Field_of_view) ;
		SIce_MY:long_name = "Multi-Year Sea Ice Concentration (%)" ;
		SIce_MY:units = "percent" ;
		SIce_MY:coordinates = "Longitude Latitude" ;
		SIce_MY:_FillValue = -999s ;
		SIce_MY:valid_range = 0, 100 ;
	short SWE(Scanline, Field_of_view) ;
		SWE:long_name = "Snow Water Equivalent (cm)" ;
		SWE:units = "cm" ;
		SWE:coordinates = "Longitude Latitude" ;
		SWE:scale_factor = 0.01 ;
		SWE:_FillValue = -999s ;
		SWE:valid_range = 0, 10000 ;
	short SWP(Scanline, Field_of_view) ;
		SWP:long_name = "Snow Water Path" ;
		SWP:units = "mm" ;
		SWP:coordinates = "Longitude Latitude" ;
		SWP:scale_factor = 0.01 ;
		SWP:_FillValue = -999s ;
		SWP:valid_range = 0, 10000 ;
	float SZ_angle(Scanline, Field_of_view) ;
		SZ_angle:long_name = "Solar Zenith Angle (-90,90) degree" ;
		SZ_angle:coordinates = "Longitude Latitude" ;
	double ScanTime_UTC(Scanline) ;
		ScanTime_UTC:long_name = "Number of seconds since 00:00:00 UTC" ;
		ScanTime_UTC:units = "seconds" ;
		ScanTime_UTC:_FillValue = -999. ;
		ScanTime_UTC:valid_range = 0., 86400. ;
	short ScanTime_dom(Scanline) ;
		ScanTime_dom:long_name = "Calendar day of the month 1-31" ;
		ScanTime_dom:units = "days" ;
		ScanTime_dom:_FillValue = -999s ;
		ScanTime_dom:valid_range = 1, 31 ;
	short ScanTime_doy(Scanline) ;
		ScanTime_doy:long_name = "julian day 1-366" ;
		ScanTime_doy:units = "days" ;
		ScanTime_doy:_FillValue = -999s ;
		ScanTime_doy:valid_range = 1, 366 ;
	short ScanTime_hour(Scanline) ;
		ScanTime_hour:long_name = "hour of the day 0-23" ;
		ScanTime_hour:units = "hours" ;
		ScanTime_hour:_FillValue = -999s ;
		ScanTime_hour:valid_range = 0, 23 ;
	short ScanTime_minute(Scanline) ;
		ScanTime_minute:long_name = "minute of the hour 0-59" ;
		ScanTime_minute:units = "minutes" ;
		ScanTime_minute:_FillValue = -999s ;
		ScanTime_minute:valid_range = 0, 59 ;
	short ScanTime_month(Scanline) ;
		ScanTime_month:long_name = "Calendar month 1-12" ;
		ScanTime_month:units = "months" ;
		ScanTime_month:_FillValue = -999s ;
		ScanTime_month:valid_range = 1, 12 ;
	short ScanTime_second(Scanline) ;
		ScanTime_second:long_name = "second of the minute 0-59" ;
		ScanTime_second:units = "seconds" ;
		ScanTime_second:_FillValue = -999s ;
		ScanTime_second:valid_range = 0, 59 ;
	short ScanTime_year(Scanline) ;
		ScanTime_year:long_name = "Calendar Year 20XX" ;
		ScanTime_year:units = "years" ;
		ScanTime_year:_FillValue = -999s ;
		ScanTime_year:valid_range = 2011, 2050 ;
	short Sfc_type(Scanline, Field_of_view) ;
		Sfc_type:description = "type of surface:0-ocean,1-sea ice,2-land,3-snow" ;
		Sfc_type:units = "1" ;
		Sfc_type:coordinates = "Longitude Latitude" ;
		Sfc_type:_FillValue = -999s ;
		Sfc_type:valid_range = 0, 3 ;
	short Snow(Scanline, Field_of_view) ;
		Snow:long_name = "Snow Cover" ;
		Snow:units = "1" ;
		Snow:coordinates = "Longitude Latitude" ;
		Snow:_FillValue = -999s ;
		Snow:valid_range = 0, 1 ;
	short SnowGS(Scanline, Field_of_view) ;
		SnowGS:long_name = "Snow Grain Size (mm)" ;
		SnowGS:units = "mm" ;
		SnowGS:coordinates = "Longitude Latitude" ;
		SnowGS:scale_factor = 0.01 ;
		SnowGS:_FillValue = -999s ;
		SnowGS:valid_range = 0, 2000 ;
	short SurfM(Scanline, Field_of_view) ;
		SurfM:long_name = "Surface Moisture" ;
		SurfM:scale_factor = 0.1 ;
		SurfM:coordinates = "Longitude Latitude" ;
	short SurfP(Scanline, Field_of_view) ;
		SurfP:long_name = "Surface Pressure (mb)" ;
		SurfP:units = "millibars" ;
		SurfP:coordinates = "Longitude Latitude" ;
		SurfP:scale_factor = 0.1 ;
		SurfP:_FillValue = -999s ;
		SurfP:valid_range = 0, 12000 ;
	short TPW(Scanline, Field_of_view) ;
		TPW:long_name = "Total Precipitable Water (mm)" ;
		TPW:units = "mm" ;
		TPW:coordinates = "Longitude Latitude" ;
		TPW:scale_factor = 0.1 ;
		TPW:_FillValue = -999s ;
		TPW:valid_range = 0, 2000 ;
	short TSkin(Scanline, Field_of_view) ;
		TSkin:long_name = "Skin Temperature (K)" ;
		TSkin:units = "Kelvin" ;
		TSkin:coordinates = "Longitude Latitude" ;
		TSkin:scale_factor = 0.01 ;
		TSkin:_FillValue = -999s ;
		TSkin:valid_range = 0, 40000 ;
	short WindDir(Scanline, Field_of_view) ;
		WindDir:long_name = "Wind Direction" ;
		WindDir:scale_factor = 0.01 ;
		WindDir:coordinates = "Longitude Latitude" ;
	short WindSp(Scanline, Field_of_view) ;
		WindSp:long_name = "Wind Speed (m/s)" ;
		WindSp:scale_factor = 0.01 ;
		WindSp:coordinates = "Longitude Latitude" ;
	short WindU(Scanline, Field_of_view) ;
		WindU:long_name = "U-direction Wind Speed (m/s)" ;
		WindU:scale_factor = 0.01 ;
		WindU:coordinates = "Longitude Latitude" ;
	short WindV(Scanline, Field_of_view) ;
		WindV:long_name = "V-direction Wind Speed (m/s)" ;
		WindV:scale_factor = 0.01 ;
		WindV:coordinates = "Longitude Latitude" ;
	short YM(Scanline, Field_of_view, Channel) ;
		YM:long_name = "Un-Corrected Channel Temperature (K)" ;
		YM:units = "Kelvin" ;
		YM:coordinates = "Longitude Latitude Freq" ;
		YM:scale_factor = 0.01 ;
		YM:_FillValue = -999s ;
		YM:valid_range = 0, 50000 ;

// global attributes:
		:missing_value = -999 ;
		:notretrievedproduct_value = -888 ;
		:noretrieval_value = -99 ;
		:cdf_version = 4. ;
		:alg_version = 4201 ;
		:dap_version = "v11r4" ;
		:Conventions = "CF-1.5" ;
		:Metadata_Conventions = "CF-1.5, Unidata Dataset Discovery v1.0" ;
		:standard_name_vocabulary = "CF Standard Name Table (version 17, 24 March 2011)" ;
		:project = "Microwave Integrated Retrieval System" ;
		:title = "MIRS IMG" ;
		:summary = "MIRS imaging products including surface emissivity, TPW, CLW, RWP, IWP, LST." ;
		:date_created = "2021-06-30T02:00:45Z" ;
		:institution = "DOC/NOAA/NESDIS/NDE > NPOESS Data Exploitation, NESDIS, NOAA, U.S. Department of Commerce" ;
		:naming_authority = "gov.noaa.nesdis.nde" ;
		:production_site = "NSOF" ;
		:production_environment = "OE" ;
		:satellite_name = "NPP" ;
		:instrument_name = "ATMS" ;
		:creator_name = "DOC/NOAA/NESDIS/STAR > MIRS TEAM, Center for Satellite Applications and Research, NESDIS, NOAA, U.S. Department of Commerce" ;
		:creator_email = "Christopher.Grassotti@noaa.gov, Quanhua.Liu@noaa.gov, Shu-yan.Liu@noaa.gov, ryan.honeyager@noaa.gov, Yong-Keun.Lee@noaa.gov " ;
		:creator_url = "http://www.star.nesdis.noaa.gov/mirs" ;
		:publisher_name = "DOC/NOAA/NESDIS/NDE > NPOESS Data Exploitation, NESDIS, NOAA, U.S. Department of Commerce" ;
		:publisher_email = "NDE_POC@noaa.gov" ;
		:publisher_url = "http://projects.osd.noaa.gov/NDE" ;
		:Metadata_Link = "NDE product-specific output file name" ;
		:references = "http://www.star.nesdis.noaa.gov/mirs/documentation.php" ;
		:history = "Tue Jul 30 17:46:22 2024: ncks -d Scanline,1,12,2 -d Field_of_view,86,94,2 NPR-MIRS-IMG_v11r4_npp_s202106300127386_e202106300128103_c202106300200370.nc output_2.nc\nCreated by MIRS Version 11.4" ;
		:processing_level = "NOAA Level 2 data" ;
		:source = "SATMS_npp_d20210630_t0127386_e0128103_b50120_c20210630015746003377_oebc_ops.h5" ;
		:time_coverage_start = "2021-06-30T01:27:38Z" ;
		:time_coverage_end = "2021-06-30T01:28:10Z" ;
		:cdm_data_type = "Swath" ;
		:geospatial_lat_units = "degrees_north" ;
		:geospatial_lon_units = "degrees_east" ;
		:geospatial_lat_resolution = "100" ;
		:geospatial_lon_resolution = "100" ;
		:geospatial_first_scanline_first_fov_lat = 62.49f ;
		:geospatial_first_scanline_first_fov_lon = 132.83f ;
		:geospatial_first_scanline_last_fov_lat = 71.26f ;
		:geospatial_first_scanline_last_fov_lon = -170.69f ;
		:geospatial_last_scanline_first_fov_lat = 63.63f ;
		:geospatial_last_scanline_first_fov_lon = 129.95f ;
		:geospatial_last_scanline_last_fov_lat = 72.94f ;
		:geospatial_last_scanline_last_fov_lon = -170.12f ;
		:total_number_retrievals = 1152 ;
		:percentage_optimal_retrievals = 0.1458333f ;
		:percentage_suboptimal_retrievals = 0.8541667f ;
		:percentage_bad_retrievals = 0.f ;
		:start_orbit_number = 50120 ;
		:end_orbit_number = 50120 ;
		:id = "ndepgsl-op-11_2021-06-30T02:00:45Z_0000001250129361_SATMS_npp_d20210630_t0127386_e0128103_b50120_c20210630015746003377_oebc_ops.h5" ;
		:NCO = "netCDF Operators version 5.0.6 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco)" ;
data:

 Atm_type =
  -999, -999, -999, -999, -999,
  -999, -999, -999, -999, -999,
  -999, -999, -999, -999, -999,
  -999, -999, -999, -999, -999,
  -999, -999, -999, -999, -999,
  -999, -999, -999, -999, -999 ;

 BT =
  22783, 22912, 24930, 25389, 25295, 24405, 23436, 23130, 22971, 22998, 
    23178, 23801, 24680, 25968, 27054, 24428, 26216, 26467, 26087, 25650, 
    25099, 24580,
  22992, 23085, 24983, 25439, 25236, 24334, 23387, 23066, 22996, 23026, 
    23185, 23865, 24766, 26000, 27006, 24436, 26241, 26340, 25957, 25657, 
    25037, 24441,
  23321, 23444, 25322, 25579, 25174, 24247, 23290, 23073, 23045, 23014, 
    23191, 23712, 24764, 26090, 27147, 24914, 26432, 26228, 25901, 25462, 
    24894, 24415,
  23199, 23336, 25346, 25579, 25090, 24108, 23318, 23088, 23025, 23041, 
    23299, 23765, 24783, 26229, 26996, 24576, 26309, 26194, 25833, 25357, 
    24878, 24287,
  22249, 22106, 25388, 25571, 24992, 23990, 23220, 23078, 23009, 22982, 
    23324, 23975, 24971, 26157, 27281, 24225, 26407, 26237, 25857, 25437, 
    24821, 24308,
  22827, 22891, 24868, 25399, 25335, 24425, 23462, 23134, 23030, 23014, 
    23121, 23723, 24459, 25950, 27069, 24455, 26191, 26468, 26123, 25730, 
    25232, 24751,
  23020, 23075, 25014, 25446, 25230, 24284, 23418, 23143, 23034, 23032, 
    23157, 23711, 24698, 26145, 27057, 24449, 26315, 26421, 26022, 25635, 
    25144, 24591,
  23347, 23414, 25153, 25552, 25165, 24200, 23399, 23129, 23060, 23089, 
    23288, 23803, 24655, 26258, 26956, 24516, 26282, 26280, 25889, 25591, 
    24983, 24420,
  23534, 23589, 25400, 25562, 25084, 24114, 23281, 23107, 23060, 23030, 
    23415, 23839, 24765, 26067, 27021, 24636, 26282, 26189, 25717, 25250, 
    24707, 24212,
  22925, 22776, 25520, 25540, 24967, 23974, 23242, 23115, 23070, 23071, 
    23293, 23953, 24891, 26166, 27121, 24662, 26313, 26044, 25612, 25224, 
    24649, 24018,
  22785, 22913, 24856, 25357, 25224, 24406, 23493, 23177, 23077, 23039, 
    23083, 23733, 24603, 25912, 26928, 24384, 26259, 26395, 26085, 25762, 
    25154, 24650,
  23083, 23212, 25050, 25421, 25187, 24293, 23460, 23139, 23046, 23043, 
    23277, 23701, 24610, 25956, 27076, 24439, 26240, 26384, 26018, 25718, 
    25080, 24463,
  23522, 23547, 25328, 25526, 25120, 24219, 23399, 23167, 23048, 23032, 
    23233, 23831, 24692, 25999, 27087, 24582, 26300, 26294, 25968, 25524, 
    24912, 24278,
  23858, 23850, 25451, 25606, 25050, 24151, 23340, 23122, 23075, 23101, 
    23232, 23764, 24926, 26166, 27335, 24755, 26276, 26145, 25769, 25431, 
    24820, 24237,
  23351, 23287, 25614, 25582, 24953, 23988, 23273, 23125, 23073, 23111, 
    23346, 23865, 24862, 26135, 27366, 24968, 26319, 26000, 25553, 25145, 
    24514, 24150,
  22691, 22869, 24796, 25340, 25240, 24398, 23500, 23176, 23101, 23078, 
    23158, 23842, 24623, 25941, 27191, 24309, 26150, 26386, 26043, 25697, 
    25245, 24645,
  23145, 23292, 25106, 25498, 25198, 24335, 23482, 23226, 23056, 23043, 
    23244, 23709, 24688, 25934, 27109, 24451, 26248, 26368, 25996, 25566, 
    25043, 24566,
  23699, 23739, 25354, 25490, 25142, 24214, 23399, 23222, 23120, 23071, 
    23290, 23844, 24789, 25938, 26644, 24535, 26147, 26292, 25906, 25503, 
    24983, 24440,
  24080, 24060, 25434, 25530, 25012, 24117, 23351, 23210, 23079, 23063, 
    23276, 23883, 24725, 25937, 27007, 24731, 26185, 26107, 25755, 25423, 
    24828, 24292,
  23592, 23565, 25572, 25530, 24914, 24021, 23295, 23171, 23101, 23070, 
    23301, 23926, 24976, 26226, 27186, 25033, 26302, 25956, 25573, 25149, 
    24618, 24037,
  22604, 22792, 24887, 25370, 25212, 24392, 23513, 23224, 23081, 23038, 
    23231, 23864, 24553, 25832, 27016, 24514, 26441, 26382, 26095, 25701, 
    25101, 24472,
  23213, 23346, 25154, 25493, 25173, 24264, 23460, 23210, 23074, 23107, 
    23115, 23794, 24659, 25703, 26934, 24801, 26347, 26313, 26041, 25570, 
    25026, 24499,
  23844, 23908, 25314, 25601, 25137, 24194, 23408, 23197, 23094, 23045, 
    23218, 23729, 24612, 26007, 26788, 24567, 26215, 26252, 25895, 25475, 
    24857, 24326,
  24154, 24118, 25323, 25525, 25001, 24094, 23339, 23146, 23156, 23086, 
    23317, 23821, 24937, 26126, 27279, 24417, 26060, 26175, 25758, 25295, 
    24848, 24252,
  23680, 23622, 25445, 25471, 24904, 24010, 23310, 23164, 23151, 23082, 
    23391, 23899, 25043, 26398, 27133, 24604, 26071, 26031, 25665, 25214, 
    24555, 24192,
  22502, 22810, 24918, 25348, 25238, 24415, 23482, 23275, 23107, 23069, 
    23266, 23749, 24689, 25772, 26984, 24746, 26381, 26425, 26097, 25654, 
    25151, 24571,
  23142, 23370, 25183, 25482, 25159, 24305, 23498, 23258, 23099, 23090, 
    23304, 23737, 24781, 25911, 27006, 24900, 26432, 26320, 25940, 25504, 
    24911, 24411,
  23857, 23971, 25382, 25533, 25138, 24234, 23450, 23222, 23155, 23120, 
    23308, 23834, 24697, 26135, 27103, 24674, 26057, 26237, 25884, 25434, 
    24908, 24446,
  24157, 24150, 25336, 25505, 25033, 24131, 23380, 23230, 23167, 23140, 
    23343, 23874, 24776, 26118, 27457, 24030, 25846, 26267, 25891, 25516, 
    24950, 24552,
  23720, 23667, 25385, 25411, 24896, 23991, 23356, 23217, 23182, 23182, 
    23423, 23942, 24912, 26132, 27319, 23902, 25670, 26015, 25648, 25242, 
    24752, 24318 ;

 CLW =
  0, 2, 0, 0, 0,
  1, 1, 0, 0, 0,
  1, 1, 0, 0, 0,
  1, 0, 0, 0, 0,
  1, 0, 0, 0, 0,
  2, 3, 0, 0, 0 ;

 ChanSel =
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1 ;

 ChiSqr =
  0.7953712, 0.59142, 0.2517513, 0.2231312, 0.2901628,
  0.83801, 0.7016711, 0.3099987, 0.3094735, 0.2798543,
  0.5025061, 0.6696218, 0.2448571, 0.2615377, 0.1434069,
  0.7199245, 0.9713045, 0.2094672, 0.3212895, 0.1872596,
  0.6445412, 0.3647941, 0.2405015, 0.3071654, 0.4628202,
  0.4326323, 0.4469193, 0.2237365, 0.4775677, 0.4854324 ;

 CldBase =
  -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888 ;

 CldThick =
  -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888 ;

 CldTop =
  -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888 ;

 Emis =
  7900, 8038, 8016, 8028, 8037, 8044, 8050, 8054, 8060, 8073, 8073, 8073, 
    8073, 8073, 8073, 8512, 8598, 8677, 8677, 8677, 8677, 8677,
  7963, 8068, 7996, 8004, 8011, 8016, 8021, 8024, 8028, 8038, 8038, 8038, 
    8038, 8038, 8038, 8435, 8493, 8571, 8571, 8571, 8571, 8571,
  7999, 8254, 8379, 8373, 8369, 8365, 8362, 8360, 8357, 8350, 8350, 8350, 
    8350, 8350, 8350, 8461, 8113, 8113, 8113, 8113, 8113, 8113,
  7962, 8214, 8414, 8402, 8393, 8386, 8379, 8374, 8370, 8355, 8355, 8355, 
    8355, 8355, 8355, 8300, 7873, 7873, 7873, 7873, 7873, 7873,
  7351, 7699, 8199, 8184, 8173, 8165, 8157, 8151, 8146, 8129, 8129, 8129, 
    8129, 8129, 8129, 8018, 7554, 7554, 7554, 7554, 7554, 7555,
  7898, 8027, 7927, 7939, 7947, 7954, 7960, 7963, 7969, 7982, 7982, 7982, 
    7982, 7982, 7982, 8485, 8512, 8594, 8594, 8594, 8594, 8594,
  8003, 8131, 8112, 8122, 8130, 8136, 8142, 8145, 8150, 8162, 8162, 8162, 
    8162, 8162, 8162, 8555, 8637, 8714, 8714, 8714, 8714, 8714,
  8096, 8287, 8291, 8286, 8282, 8279, 8277, 8274, 8272, 8267, 8267, 8267, 
    8267, 8267, 8267, 8316, 8066, 8066, 8066, 8066, 8066, 8066,
  8140, 8362, 8497, 8483, 8474, 8467, 8460, 8455, 8450, 8435, 8435, 8435, 
    8435, 8435, 8435, 8352, 7930, 7930, 7930, 7930, 7930, 7930,
  7763, 8105, 8563, 8542, 8528, 8517, 8506, 8498, 8490, 8467, 8467, 8467, 
    8467, 8467, 8467, 8325, 7682, 7682, 7682, 7682, 7682, 7682,
  7887, 8009, 7952, 7963, 7971, 7977, 7983, 7986, 7991, 8003, 8003, 8003, 
    8003, 8003, 8003, 8438, 8510, 8591, 8591, 8591, 8591, 8591,
  8099, 8224, 8247, 8257, 8264, 8270, 8275, 8278, 8283, 8294, 8294, 8294, 
    8294, 8294, 8294, 8619, 8726, 8799, 8799, 8799, 8799, 8799,
  8227, 8432, 8531, 8521, 8514, 8509, 8504, 8500, 8496, 8485, 8485, 8485, 
    8485, 8485, 8485, 8426, 8109, 8109, 8109, 8109, 8109, 8109,
  8360, 8576, 8694, 8677, 8665, 8656, 8647, 8641, 8635, 8616, 8616, 8616, 
    8616, 8616, 8616, 8494, 7976, 7976, 7976, 7976, 7976, 7976,
  7969, 8301, 8708, 8687, 8673, 8662, 8651, 8644, 8636, 8613, 8613, 8613, 
    8613, 8613, 8613, 8502, 7840, 7839, 7839, 7839, 7840, 7840,
  7890, 8017, 7942, 7953, 7962, 7968, 7974, 7977, 7983, 7996, 7996, 7996, 
    7996, 7996, 7996, 8465, 8517, 8598, 8598, 8598, 8598, 8598,
  8123, 8254, 8310, 8320, 8328, 8333, 8339, 8342, 8347, 8358, 8358, 8358, 
    8358, 8358, 8358, 8658, 8784, 8856, 8856, 8856, 8856, 8856,
  8341, 8534, 8596, 8582, 8573, 8565, 8558, 8553, 8548, 8533, 8533, 8533, 
    8533, 8533, 8533, 8434, 8021, 8021, 8021, 8021, 8021, 8021,
  8579, 8781, 8864, 8845, 8831, 8821, 8811, 8804, 8796, 8775, 8775, 8775, 
    8775, 8775, 8775, 8620, 8049, 8049, 8049, 8049, 8049, 8049,
  8177, 8492, 8840, 8819, 8805, 8794, 8783, 8775, 8768, 8745, 8745, 8745, 
    8745, 8745, 8745, 8643, 7969, 7969, 7969, 7969, 7969, 7969,
  7773, 7931, 7968, 7982, 7993, 8001, 8009, 8013, 8020, 8036, 8036, 8036, 
    8036, 8036, 8036, 8484, 8625, 8708, 8708, 8708, 8708, 8708,
  8087, 8316, 8371, 8372, 8372, 8372, 8372, 8371, 8371, 8371, 8371, 8371, 
    8371, 8371, 8371, 8550, 8369, 8369, 8369, 8369, 8369, 8369,
  8361, 8528, 8523, 8512, 8504, 8498, 8492, 8488, 8483, 8471, 8471, 8471, 
    8471, 8471, 8471, 8389, 8047, 8047, 8047, 8047, 8047, 8047,
  8572, 8705, 8646, 8630, 8618, 8609, 8600, 8594, 8588, 8569, 8569, 8569, 
    8569, 8569, 8569, 8377, 7939, 7939, 7939, 7939, 7939, 7939,
  8341, 8582, 8778, 8757, 8742, 8731, 8719, 8711, 8704, 8680, 8680, 8680, 
    8680, 8680, 8680, 8501, 7873, 7873, 7873, 7873, 7873, 7873,
  7735, 7906, 7915, 7931, 7943, 7952, 7960, 7965, 7972, 7990, 7990, 7990, 
    7990, 7990, 7990, 8514, 8625, 8711, 8711, 8711, 8711, 8711,
  8038, 8195, 8277, 8290, 8299, 8306, 8313, 8317, 8323, 8338, 8338, 8338, 
    8338, 8338, 8338, 8696, 8838, 8912, 8912, 8912, 8912, 8912,
  8463, 8662, 8709, 8695, 8685, 8677, 8670, 8664, 8659, 8643, 8643, 8643, 
    8643, 8643, 8643, 8574, 8101, 8101, 8101, 8101, 8101, 8102,
  8699, 8838, 8796, 8776, 8762, 8751, 8741, 8733, 8726, 8704, 8704, 8704, 
    8704, 8704, 8704, 8478, 7953, 7953, 7953, 7953, 7953, 7953,
  8548, 8757, 8934, 8904, 8884, 8868, 8852, 8842, 8831, 8798, 8798, 8798, 
    8798, 8798, 8798, 8444, 7684, 7684, 7684, 7684, 7684, 7684 ;

 Freq = 23.8, 31.4, 50.3, 51.76, 52.8, 53.596, 54.4, 54.94, 55.5, 57.29, 
    57.29, 57.29, 57.29, 57.29, 57.29, 88.2, 165.5, 183.31, 183.31, 183.31, 
    183.31, 183.31 ;

 GWP =
  _, _, _, _, _,
  _, _, _, _, _,
  _, _, _, _, _,
  _, _, _, _, _,
  _, _, _, _, _,
  _, _, _, _, _ ;

 IWP =
  _, _, _, _, _,
  _, _, _, _, _,
  _, _, _, _, _,
  _, _, _, _, _,
  _, _, _, _, _,
  _, _, _, _, _ ;

 LWP =
  -998, -998, -998, -998, -998,
  -998, -998, -998, -998, -998,
  -998, -998, -998, -998, -998,
  -998, -998, -998, -998, -998,
  -998, -998, -998, -998, -998,
  -998, -998, -998, -998, -998 ;

 LZ_angle =
  50.16999, 53.05, 56.09, 59.2, 62.46,
  50.15999, 53.08001, 56.07, 59.21998, 62.46,
  50.14001, 53.08001, 56.08001, 59.2, 62.48999,
  50.15999, 53.06001, 56.09999, 59.18999, 62.46998,
  50.16999, 53.07, 56.08001, 59.21, 62.46,
  50.14001, 53.09001, 56.07, 59.21998, 62.46998 ;

 Latitude =
  71.45, 71.51, 71.54, 71.53, 71.47,
  71.76, 71.82, 71.85, 71.84, 71.78,
  72.07, 72.13, 72.16, 72.15, 72.08,
  72.38, 72.44, 72.47, 72.46, 72.39,
  72.69, 72.75, 72.78, 72.77, 72.7,
  73, 73.06, 73.09, 73.08, 73.01 ;

 Longitude =
  176.67, 178.83, -178.67, -175.83, -172.53,
  176.55, 178.78, -178.72, -175.8, -172.46,
  176.43, 178.7, -178.75, -175.81, -172.36,
  176.32, 178.6, -178.76, -175.8, -172.31,
  176.21, 178.53, -178.82, -175.76, -172.25,
  176.07, 178.46, -178.86, -175.74, -172.14 ;

 Orb_mode = 0, 0, 0, 0, 0, 0 ;

 Polo = 2, 2, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 2, 3, 3, 3, 3, 3, 3 ;

 PrecipType =
  -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888 ;

 Prob_SF =
  _, _, _, _, _,
  _, _, _, _, _,
  _, _, _, _, _,
  _, _, _, _, _,
  _, _, _, _, _,
  _, _, _, _, _ ;

 Qc =
  0, 0, 0, 4096,
  0, 0, 32, 4096,
  1, 0, 144, 0,
  1, 0, 144, 0,
  1, 0, 144, 0,
  0, 0, 0, 4096,
  0, 0, 0, 4096,
  1, 0, 144, 0,
  0, 0, 128, 0,
  1, 0, 144, 0,
  0, 0, 0, 4096,
  0, 0, 0, 4096,
  1, 0, 144, 0,
  1, 0, 144, 0,
  1, 0, 144, 0,
  0, 0, 0, 4096,
  0, 0, 0, 4096,
  1, 0, 144, 0,
  1, 0, 148, 0,
  1, 0, 156, 0,
  1, 0, 20, 4096,
  1, 0, 144, 0,
  1, 0, 144, 0,
  1, 0, 144, 0,
  1, 0, 144, 0,
  0, 0, 32, 4096,
  0, 0, 32, 4096,
  1, 0, 144, 0,
  1, 0, 144, 0,
  1, 0, 144, 0 ;

 RAzi_angle =
  -95.24, -93.2, -90.83, -88.14, -85.01,
  -95.3, -93.19, -90.81, -88.04, -84.86,
  -95.35, -93.19, -90.76, -87.97, -84.69,
  -95.4, -93.22, -90.71, -87.89, -84.56,
  -95.44, -93.22, -90.69, -87.77, -84.42,
  -95.51, -93.22, -90.66, -87.68, -84.24 ;

 RFlag =
  -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888 ;

 RR =
  _, _, _, _, _,
  _, _, _, _, _,
  _, _, _, _, _,
  _, _, _, _, _,
  _, _, _, _, _,
  _, _, _, _, _ ;

 RWP =
  _, _, _, _, _,
  _, _, _, _, _,
  _, _, _, _, _,
  _, _, _, _, _,
  _, _, _, _, _,
  _, _, _, _, _ ;

 SFR =
  _, _, _, _, _,
  _, _, _, _, _,
  _, _, _, _, _,
  _, _, _, _, _,
  _, _, _, _, _,
  _, _, _, _, _ ;

 SIce =
  76, 76, 80, 80, 66,
  76, 78, 80, 82, 78,
  76, 82, 84, 88, 82,
  76, 82, 88, 94, 88,
  74, 82, 86, 90, 88,
  74, 82, 90, 94, 92 ;

 SIce_FY =
  76, 76, 80, 80, 66,
  76, 78, 80, 82, 78,
  76, 82, 84, 88, 82,
  76, 82, 88, 94, 88,
  74, 82, 86, 90, 88,
  74, 82, 90, 94, 92 ;

 SIce_MY =
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0,
  0, 0, 0, 0, 0 ;

 SWE =
  _, _, _, _, _,
  _, _, _, _, _,
  _, _, _, _, _,
  _, _, _, _, _,
  _, _, _, _, _,
  _, _, _, _, _ ;

 SWP =
  _, _, _, _, _,
  _, _, _, _, _,
  _, _, _, _, _,
  _, _, _, _, _,
  _, _, _, _, _,
  _, _, _, _, _ ;

 SZ_angle =
  49.34, 49.66, 50.03, 50.46, 50.97,
  49.62, 49.94, 50.3, 50.73, 51.24,
  49.9, 50.22, 50.58, 51, 51.51,
  50.18, 50.49, 50.86, 51.27, 51.78,
  50.46, 50.77, 51.13, 51.55, 52.05,
  50.74, 51.05, 51.4, 51.82, 52.32 ;

 ScanTime_UTC = 5261.00048828125, 5266.00048828125, 5272.00048828125, 
    5277.00048828125, 5282.00048828125, 5288.00048828125 ;

 ScanTime_dom = 30, 30, 30, 30, 30, 30 ;

 ScanTime_doy = 181, 181, 181, 181, 181, 181 ;

 ScanTime_hour = 1, 1, 1, 1, 1, 1 ;

 ScanTime_minute = 27, 27, 27, 27, 28, 28 ;

 ScanTime_month = 6, 6, 6, 6, 6, 6 ;

 ScanTime_second = 41, 46, 52, 57, 2, 8 ;

 ScanTime_year = 2021, 2021, 2021, 2021, 2021, 2021 ;

 Sfc_type =
  1, 1, 1, 1, 1,
  1, 1, 1, 1, 1,
  1, 1, 1, 1, 1,
  1, 1, 1, 1, 1,
  1, 1, 1, 1, 1,
  1, 1, 1, 1, 1 ;

 Snow =
  _, _, _, _, _,
  _, _, _, _, _,
  _, _, _, _, _,
  _, _, _, _, _,
  _, _, _, _, _,
  _, _, _, _, _ ;

 SnowGS =
  _, _, _, _, _,
  _, _, _, _, _,
  _, _, _, _, _,
  _, _, _, _, _,
  _, _, _, _, _,
  _, _, _, _, _ ;

 SurfM =
  -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888 ;

 SurfP =
  10084, 10084, 9930, 9930, 9930,
  10084, 10084, 9930, 9930, 9930,
  10084, 10084, 9930, 9930, 9930,
  10084, 10084, 9930, 9930, 9930,
  10084, 9930, 9930, 9930, 9930,
  10084, 10084, 9930, 9930, 9930 ;

 TPW =
  96, 104, 134, 128, 130,
  100, 101, 123, 124, 131,
  103, 94, 125, 130, 132,
  99, 94, 115, 129, 138,
  116, 123, 119, 110, 113,
  104, 106, 111, 99, 103 ;

 TSkin =
  27765, 27612, 27572, 27487, 27762,
  27740, 27634, 27429, 27474, 27567,
  27662, 27494, 27256, 27280, 27575,
  27628, 27562, 27275, 26996, 27279,
  27697, 27310, 27381, 27248, 27204,
  27713, 27563, 27188, 27092, 26923 ;

 WindDir =
  -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888 ;

 WindSp =
  -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888 ;

 WindU =
  -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888 ;

 WindV =
  -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888,
  -888, -888, -888, -888, -888 ;

 YM =
  23075, 23066, 25066, 25344, 25162, 24317, 23365, 23011, 22865, 22945, 
    23118, 23752, 24605, 25872, 26984, 24490, 26046, 26310, 25960, 25533, 
    24987, 24516,
  23295, 23256, 25067, 25355, 25091, 24245, 23311, 22944, 22889, 22972, 
    23122, 23813, 24689, 25904, 26932, 24464, 26065, 26179, 25831, 25541, 
    24924, 24377,
  23616, 23622, 25341, 25449, 25017, 24156, 23210, 22947, 22936, 22958, 
    23125, 23657, 24682, 25989, 27074, 24882, 26239, 26057, 25769, 25342, 
    24778, 24351,
  23539, 23574, 25298, 25396, 24923, 24008, 23235, 22960, 22913, 22985, 
    23231, 23707, 24697, 26122, 26921, 24479, 26097, 26015, 25694, 25237, 
    24759, 24218,
  22665, 22444, 25263, 25351, 24817, 23885, 23131, 22948, 22897, 22925, 
    23257, 23913, 24880, 26048, 27204, 24054, 26184, 26051, 25715, 25312, 
    24697, 24232,
  23119, 23045, 25004, 25354, 25202, 24337, 23391, 23015, 22924, 22961, 
    23061, 23674, 24384, 25854, 26998, 24517, 26021, 26310, 25997, 25613, 
    25120, 24687,
  23323, 23246, 25098, 25362, 25085, 24195, 23343, 23021, 22927, 22978, 
    23094, 23659, 24621, 26050, 26984, 24477, 26139, 26260, 25895, 25520, 
    25031, 24527,
  23642, 23592, 25172, 25422, 25008, 24109, 23319, 23004, 22951, 23033, 
    23222, 23748, 24573, 26157, 26882, 24484, 26090, 26110, 25757, 25471, 
    24867, 24355,
  23874, 23827, 25352, 25379, 24917, 24014, 23198, 22979, 22948, 22974, 
    23348, 23781, 24679, 25960, 26946, 24539, 26071, 26010, 25578, 25130, 
    24588, 24142,
  23341, 23114, 25395, 25320, 24792, 23869, 23153, 22985, 22958, 23014, 
    23226, 23891, 24800, 26057, 27045, 24491, 26090, 25859, 25469, 25099, 
    24525, 23942,
  23077, 23067, 24992, 25312, 25091, 24318, 23422, 23058, 22971, 22986, 
    23023, 23684, 24528, 25816, 26857, 24446, 26088, 26238, 25959, 25645, 
    25042, 24586,
  23386, 23383, 25134, 25337, 25042, 24204, 23384, 23017, 22939, 22989, 
    23214, 23649, 24533, 25860, 27003, 24467, 26064, 26224, 25891, 25601, 
    24967, 24399,
  23817, 23725, 25347, 25396, 24963, 24128, 23319, 23041, 22939, 22976, 
    23167, 23776, 24610, 25898, 27013, 24550, 26107, 26124, 25835, 25404, 
    24796, 24213,
  24198, 24088, 25403, 25423, 24883, 24051, 23257, 22994, 22963, 23045, 
    23164, 23706, 24840, 26059, 27260, 24658, 26065, 25966, 25629, 25311, 
    24701, 24167,
  23767, 23625, 25489, 25362, 24778, 23883, 23184, 22995, 22961, 23054, 
    23279, 23803, 24771, 26026, 27290, 24797, 26096, 25815, 25410, 25020, 
    24390, 24074,
  22983, 23023, 24932, 25295, 25107, 24310, 23429, 23057, 22995, 23025, 
    23098, 23793, 24548, 25845, 27121, 24371, 25979, 26229, 25917, 25580, 
    25133, 24581,
  23448, 23463, 25190, 25414, 25053, 24246, 23406, 23104, 22949, 22989, 
    23181, 23657, 24611, 25839, 27035, 24479, 26072, 26207, 25869, 25450, 
    24930, 24502,
  23994, 23917, 25373, 25360, 24985, 24123, 23319, 23096, 23011, 23015, 
    23224, 23789, 24707, 25837, 26571, 24503, 25954, 26122, 25774, 25383, 
    24867, 24375,
  24420, 24298, 25386, 25347, 24845, 24017, 23268, 23082, 22968, 23007, 
    23208, 23825, 24639, 25829, 26932, 24634, 25974, 25928, 25616, 25303, 
    24709, 24222,
  24008, 23903, 25447, 25310, 24739, 23916, 23206, 23041, 22989, 23013, 
    23234, 23864, 24885, 26118, 27110, 24862, 26079, 25770, 25430, 25024, 
    24494, 23962,
  22896, 22946, 25023, 25325, 25079, 24304, 23442, 23105, 22975, 22985, 
    23171, 23815, 24478, 25737, 26945, 24576, 26270, 26225, 25969, 25584, 
    24989, 24408,
  23516, 23517, 25238, 25409, 25028, 24175, 23384, 23088, 22967, 23054, 
    23052, 23742, 24582, 25607, 26860, 24829, 26171, 26153, 25914, 25454, 
    24913, 24435,
  24139, 24086, 25333, 25471, 24980, 24103, 23328, 23071, 22985, 22989, 
    23152, 23674, 24530, 25906, 26715, 24535, 26022, 26082, 25763, 25355, 
    24741, 24262,
  24494, 24356, 25275, 25342, 24834, 23994, 23256, 23018, 23044, 23030, 
    23249, 23763, 24851, 26019, 27204, 24320, 25848, 25996, 25619, 25175, 
    24729, 24182,
  24096, 23960, 25320, 25251, 24729, 23905, 23221, 23034, 23039, 23025, 
    23324, 23837, 24952, 26289, 27057, 24433, 25848, 25845, 25522, 25089, 
    24431, 24116,
  22794, 22964, 25054, 25303, 25105, 24327, 23411, 23156, 23001, 23016, 
    23206, 23700, 24614, 25676, 26913, 24808, 26210, 26268, 25971, 25537, 
    25039, 24507,
  23445, 23541, 25267, 25398, 25014, 24216, 23422, 23136, 22992, 23037, 
    23241, 23685, 24704, 25816, 26932, 24928, 26256, 26160, 25813, 25388, 
    24798, 24347,
  24152, 24149, 25401, 25403, 24981, 24143, 23370, 23096, 23046, 23064, 
    23242, 23779, 24615, 26034, 27029, 24642, 25864, 26067, 25751, 25314, 
    24792, 24381,
  24497, 24388, 25288, 25322, 24866, 24031, 23297, 23102, 23055, 23084, 
    23276, 23816, 24690, 26010, 27382, 23933, 25634, 26088, 25751, 25396, 
    24831, 24482,
  24136, 24005, 25260, 25191, 24721, 23886, 23267, 23087, 23070, 23125, 
    23356, 23880, 24821, 26023, 27243, 23731, 25447, 25829, 25505, 25117, 
    24628, 24242 ;
}
